XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180�Em�qǹ㢮
Xq�$��V�)�Qj�C՜�<ZQ�3��d����"�6���=h���o��
���jO}=؁�M�s�p��95q��
fl�Q��,G���\x{�9]���@u�A&N��D1��4�"�EH�������h0y�^�l�UAZ�=Z$��-�%i�1�)�ƔY#2 �^H���*p�t'F���q�d0V+�z���GT��s[dP�F3�Ф�#j��t.��f ����TE�a����YB�Z�<�Q@����ػ�@�?�W�ׅ9 !d��J�ȗ�7�d���SЛ�^8�A��M2s54���/eM����ҶH�i	@u�Ҽ��C�O>�;[��&a8Hl��L`C��`0Е=���Eֿ��XlxV61EB     400     130�����UK���Z����3=U$|���3�̽bG����c�B
^�Ìԁ����-����o�=σn�0��I}��|��-K�${�Eo�Wf<K��v�U���F��fV��U�����T�y�P�@h�]����4��YxGǤ�y����qR���gGp�;�L�P&�R�Nd4�bcr#-�ی�_&���W	��@a���NA|e�����:�,�xf;����eh�a���R�pNr�Cc3��\.�P�FJr[
l:���^c�u�Ļ/�`�[�(��Ѽ�W�SX�%�iB*�XlxV61EB     400     190:�~�rT��AY��VA�=�.<N����r�a�\S�*	s�IJ=�-�愦-�'9q�ƴ|��y�y�
~����ZwĩMZ�*������Q:p;�z�'��"r�.�b�v�/;�lyZ�yTe��	�Kq
%¾?�ٔ�*[q�8���W�zCL]��@� �R���ݝe�S� �ۚ�h�q�m��4����zA�i����'��m��Y�%�ׁ1DP�P0�Oڽ ��!��D�hrǇZ�W�w
�"Y̎�ɜq�����R\e��'�|��P;$A[A��T"t�����pj�]N�9��κ���;BN��{1Bul��s����౬$��w߂�� ���v���O>|x�	�]� �k�E������9��g*T�� U�%mDT�q�#V�ܜ9�Y}TXlxV61EB     400     1308�l|��M�EI�j���m�֛)�Y�9���&4pe��)8�˼��vЧfVN�!����I����4�rE�]�@2�:_����	���k���.��Maw�x�n7Fe(�O�C���C�z�BF|���ƚ�Z�4�����c�p~�.q�O_\yR1���T{ou��r*�lGf{��+�.�j�!��3�ٍ���#s�PAlq �B&�mըܲ����:�Qkج�iN,n ��F���c�a"�t/6q�z�O��S+�<ﾺ�oJZTVz��s���j�t���muxkk��L�pJ���XlxV61EB     400     110��Bv?2���a�)���}�U&��\�L��vKjX����.�!W�0��� |�1��x�q��0�DL31�����<����EuWzb�Ou�I��,.�ټ{��(���eq����j�D: 'hԡn �Z��Bq������R7��1���zJ�M|ܢ�Q͝�8�,�b�@&D��W�3�pč���N��2����fؘZ��{koݫl�'��z�,��ǩ�d��Z�4��-x�gE+����PG[�g���v��{�)]���:tXlxV61EB     400     190n������7Y�e�w��EQP6ez�]݄��o��b�@�r���^����5�2��m�I��p�8�fg\u��Z�<���`��,w��Nq��� _ �E���UGH����ƾ���Ft�sJ� �I\\M�,�=׭e��ơϕ
��$��_xp���6���dn�}
���^D��M�� �dO��ɕʊ�m�^��߻�U	F�B�z��h�(v\Ÿ�t�C�x|=9zm�q�z���%�o�M�O:x3���� \H�Y��:w� h֩�D��Y?f��p��:�b�xh�%q-����T��8&4��T.�3ht�YC|�SN<��:Q�g�6��dt�H��f̿j�Y�llż̦�D��m}n�!��RzqU��ew�}�`�80�=��CXlxV61EB     400     160�&�l�[o��Z�j0� �Nz�!�t�z=��๫���;�p�MU�����������B�);�O:�C��Db7�9�Vʻv}�Ԁ���<3e�G�G��wv����dH���+D��@��8+x�o�N�9VϜh�sq'�k�m9�B&�ַ���[:�.��´c�ҟad�~ճTiNRc����X���yl����3�w�E� Z�&���bF��Y>��ړ�w2�J���z��A�Z��r�ƄS��Dg52���܏�I�o}�g4,cn]Nh��6qC�AJ^9L2�_�6�G����Cc�+e�ضRoJcP�7f�1�Ϯûj��ܽlגK�:�]Mv��XlxV61EB     400     1c0�zf��3�x��x��0���z#�;�K��4��>-���~��G$���u�ڈc\��`D9|-�q��%�����U�S�����V�[�����zt�,��ļ�As��(�y��j�XI��6P����e��˼����⊝��%��D0˹38wK�&��I�C9/
�4^Im�d�+*��i�
�y�ƀt�No� ����{���!Y7���;�e]x���
)�a���͛#���jȘ� �+�J�޹�s]l�j���#��Yeh�Y�8X�< ��	�'
4�`��ͬ��K�}��+�A2"ƚ3�YW�@(b�Xԅ��*@:O�*�c4��&hD
�ͫ#a�m�~>ZrT}B���b�A�<�����/_�W{��ŝCBM�Vɳ�B�r����9E'Ft'R�3!> �b�[Ȣ�ϫ��Pm��`T[�8.����x�X/|XlxV61EB     400     1c0ڍpL�V'7�|Q,t�/�e�7a{��9�?>43U(W�k鮣����!v�s��~*�|���d��+�;^���L~ ���X	q�cϷ��դ�Ʋ����q����y3nW <����y���T�E8��8M���R��u�D��9Ě@���D�>���[:�w�$<�@�>O�|M�3��c�����n��.�����t�6炛(�q,��@�������, O��pk�E�
�=�#�������Q��*ř)G������S(k�c#�sޘP%UH�U�Ⱦ��B��E���<�v.f
����P�ݖ	��vO��[��d3?;oe2�)ݦu�i&w=�>~ �vZ�V7}���I{��h��L����;:�qB�f�G��hk~=�5�E�-�%M����g(��P'�'%m�M~����g�A4Sx����4	�3�XlxV61EB      ef      a0p��v�Qw�<I�?9�|z�_�-j����8$n�h���Mz����w5Orz�>�2�@�Ceӓ��҉6[|�*� $�u�8ߗ:1K����� ̻؎�i��@x^�4�Hӧ�;��׊&RxĿ���?�Ʉ���c�o�I�5}[��A*PG��/����