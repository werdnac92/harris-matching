XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160��Te}���i~�?����ak���e+�A^L%l�;qEA|J���з�x��W���,��x��i'�ؘ&�ү��6Xj�;��s�XM�b�*���aN�,����igp��
�;�j��:��*LKkxԜ~��s�Tc�Vs�.�c�e��T(C��/r�2o5Jwh�d����d5.
�<���[p$pңUk���H{�������ui�$1B脕��'ݲu1ʪ�+!]�q��d���s�(�.��'m:2���+�Z���@�e5��]-ڐv��/�&od���'6�Zd�����Z<��TI�!x��o�a���0�.WT���a[�ϕ"*�XlxV61EB     400     160��'�uEN��W'I��ܟu��Ix�Ӵ�O�.���v�|Ӯ���z�srB<F�c�7s�FI8���=����oД%U�Q����W�k��N���u�-%0*��믱;���pX�E���:9�}Ձ��/�ޓ����	���'n{�'��?�k������u�S��)��BO���/��*.i��h�'a��+�7�l��9#YC�~���V0;�����$�9�*)���>t���ݣ�I�w�y���BL�YX���� p��k�\���Ux-/�-�����q��3<�u�z���zH��8���6�<alW7��7���cd��ChT>dXlxV61EB     400      e0Z{g{$c��M�}�P�	�*�~�7�6��Q�^�L�!0܎�XN���T�!�����A0�{�k�jz���8?-�@h�>ŷ�<���|Sf����&�ɹYqw�+A˟b"���2D�*O�g�G�6:�L�H]	�ypȢA�xS�1;3Mv��:f$?�͛����y�}j0�Fh��NSc/�F�l (��7Rf����y�p�|�NE�\7/�/XlxV61EB     400     160�9����ce q��n!@��'��X���+�y�'���L� ��`����ӣ�Pu���ڰΐY��u�ړy�Sm:uy������-9�����e`�?���wC�۩xĨ ���g��/�[�d����,�0ֲ5�I����p�Aw
>G�=�H�⍪]z!�fW�e4�i"�!�	���x�^�v��,�kr�(��I�C�p�uϕ����,���7�7kE����؏��50�y9a���2�),=��p�����7���v�~ �頍�ٻvu�-y]6?iгb�cc��e~8���;�'��˧ń^���wk̻�-���6��r��_!cB��B��p�s߭��F[4�EXlxV61EB     400     150^�\N]vX( X�U��W��zr���	;�2?��i/�Bfoz�đ�`I�����X;�0��Sz]�Ô��d�-�sڱud�@��"��C�Q����
���Mܨd!^�Ӽ�`El���п?�_B?���%����� H�/���m��;�M�T�*E�5l�i��-����.��B��Z��p=e��.�A�z��p7�Z/o��<F��`ҁ����9y�����q}d"�I.�� ?b1���$H��ل���������
A3�L�lLI��[����+�����lr�5�~"�������,�B�Sn�S.tǋ��1�~zKrU����k�/�XlxV61EB     400     170�9�Ç���'�'N� ��[��u�����"�!'�X`8�;�����?�%m��eU���n��HTۢW����~�R� ��B]��q���dr�!��M��,l>r�%���\ml����b�(v����Q4�Z�p ����R�
�!�wY5cc?��l�sz5�3�o�/��x��5�y�K�C~���d�]����)������5D�@�;�7��tR�y8.B��/ Ʊ�6����?���ؚ �2�J!����N�en�(\g�Ʌi��"���bi�W� ��+D�sfH.m��^e{.����4�\*\� ��X��ZyT�Y=~k��JD�1N0A���#�i��t�ɧD�3)=XlxV61EB     400      b0�M�𔮃�+�)G�[��{�~�j��}ۓT;�H��R�'r!`�	6)Xw�( ,���dKL��}}�d��I��+SU��I���E��J�5�Vbg�U�A��NSZf�3ʅ�g@$���՗��+�b���f�	C�/�4:�\�O宼�7����ihOM�}���̪%G�XlxV61EB     400      c030�t/��c�:���+���6��`ߍ/�T���\rT=��R#�zD�'heaUw~��t�>¬~���T;�����Þ@�I�?%i<Ƥ�foU��rtXc��k9i�:Y�f4�ؖ�l�X�޾3ʡ8w0ܔ�FsI���q��h����(�^pw&�4�dvr#Q�����0�$���Ev��cGO�
��-��e��XlxV61EB     400      c030�t/��c�:���+��,[\��E��M���$�ݨy��__��V ��2��H��fv��v�Z��E��
O(����Yx4J��
g?��~j��,t���|��l��� �M
��5�c8�P���?�����&�)ĸ���� |{�^f��#�4�a-�p����QH��DL��I�+[��XlxV61EB     400      c00�g��s�o���|E]�0l�5=��3q�ý�B{G�=*1n$6���㩋	£fW�+Ǩ�Ci��(|�QU��(>�~Ar鑴�,����4`�L'��'�_���2��Cr�s&}�:�A������!Ǆb��+r���P�,t&�!������Y1�<V�[}'��c 2Һ�	�~�`P�XlxV61EB     400      c0�.�O��ti���b�.�q��[O��R$��]_�a>�|���@~��ϐ���/� ���`�%[Y����]�T-������8;i������^�>�Ƚؕ�"�],���*nAl���I�=��f�������[*�;s�l�6!į��2�B��p�Z}&aկ�04:Ο�~!�h��}�h����9�T��
XlxV61EB     400     1a0d��Lʨ��~`愆�]��9��+�����X}Ѻ��������<:\��\i�0�`�]�kv�n�v�J�@��n"����t�B�x1 �p?�L;�E�ҡ�l46I��-`7�N<�:-��)%�A�ovs����J���3�e�%� �_��]���%I�(M��B�h׮L�jݝX�?��ӊ}v6�nҙ*�S݅�A9nwT�d�<� @0K�HR����hV��V��Z�&n��+¾j0	���4��F抃3sX�.�-٨����� �x�@l��K�g����;�*;ꁸ�s8��]�˗� �DRXj�EwT��$��ԄY}�O#7�\��>�V�����v�{*�:��x�z#j	ӆ�8Jے��OmG�"�l��Jeȥ;Re��L��a��h���8XlxV61EB     400     150a���uUV<&fD7h·x����81��ƾO ��c(��L{�9g�A1�`[պ{����!|'�6��[��)P��-Y	��������q��r����.(pI D"N?k�]��+�0�m�~��]r`#�8.���q��1����߆\�&�y��?z�'*�nP�m��������k�P���$(*�[���%�
�ɤ�����v����V�URr�Ȟ��D��h�5Q ӳ�M�p��o��_����z�sV�׉�D�f��H��a/�["3Y7����l�^��Ԃb��N�Z��3��J8f������b9x{�cF�:U�ԩ���[XlxV61EB     400     140q�oJ+F ,�%��(�o|�؞�-������#��mz%�S�����N�����9N����C������^�<ή�ū�<^�q@6رj'8�9�������\��*�]@�1��PI9 �g��T�d���#��'q�	M=�gR��~H��Ctr�6��s�-���/8K�9�~�����/�WY�����q��"�1��+>XF��Ez�bJ��P>x�Z�"��"�����r�}��s_�o��Q&��i�zk2<3�_�b������:#��t*�ߢL�����B�]�=����׏:�}����C�a��d�Q��˖��/�<�XlxV61EB     400     130#;��k�n0ΌW���p\=~���� ۢ����3=�������H@���G爜B�O�ܢL���b����AVE�Q��bb����1Ĳ˂K�2gS~I;��.\e-@��O�b���o,Hv�V ^� �<���5�Ծr �D��L�)(�F��yكnzA`G'�����j4�n�Tπ@D����)�W�m����x��L��5J��c"/�J��+YLZB�e�VbH��;{ts����0��*n���=�+x�<Jj�Q`�싱�T����5)��Iq��f��[���xXK�R�XlxV61EB      4b      40ʒ:�ɖ�`e�%L�Zl��Pi�2H�J<9q8~��������X(P����rǅ�H