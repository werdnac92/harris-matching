XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150�I�;g�t�?g�E�cՒܮ4$͊y���햕�b�J��\�{+�2�b��e��/��(H�6`EP��(�����(�3��]�\�1t���e�Q6����E�U1S	�d~I��P��3���X72�_�?G'��
��n.0�� }m�4������bn$���F79(���M[o��L	�`��c�{0�/��3�Iz��H�����I�k^av���:�BT ���Н�N�t�Jm#4+#�Y���Oe����Ǐ�[���-��ҁ#|jR�vփ:�,R�\B�����F
�
�V{1�MG� �ѧ���g��W?��iv�8��XlxV61EB     400     140�q���už���hk ��?Y5���n)�(�<���gT��>06��`��]S�3����)�����k�2q��(����:�f�Dp�Y����h�I����"���9}˕�%��P̳������X,C�U�.���0�Q}x5����mv�j`.c�1ܺz��n���W�E�.�}Y��m���KT�I��7rnn-��vP^�V1�<=��\WN-��%T��(�����V�?a}��P1/��f�2���o7ʒ�n��ZO�e��Z�B���W�\������Ȼ!���HY�-D�E*�*��	J�XlxV61EB     289      c0-SS¹!��b�Ʉ��F����`����O�M]GE�������F0�{�\��1zJ�X��y�s�yvyj�#����L�H�+(;~�** �w����hT����S4�t9��z���q�����3[;.:'RϮp�`��D^Y��`K���pP.	���(;�6��2��O�;�y�Y#C�U��1Ùr�����