XlxV61EB     400     130D9ɛ���l�k����ͦSx�%�܄A���Gνu�Ƈ���U��8��{�מ��^Ls�&�| ����������|CJL����O ����E��Z:��; ��H�9�8��>cR���d�$(0Xe�9S� ���
Fq5��kx2rx�oS��Ѯ�XCm��A��T��0PRSuÅ�7�T(a�3 *�wʬ�j#��/������	��e��wUBm�jv��A�DŴ�;Ġ�o��;�G����`I�S����e�X�CW8�o��vp\,�L>ʭ��mb�%�C-"�����XlxV61EB     400     1d0Bf'����5�L�a 0y_ ����v�����gEΪ�}>x#ݢ3�X:Q(�Ks	�sq�.\��������;���ݐ_�/�ͺ(oe�%��>�X2�Y��ѿMi�0��5M�.wC����f�Bo3T�TK.��ń��`�-u^fZ'�=Ec�Z��b�'��q�YAI~�S�UL9>VR(#6C_�̛!�[^˷��1�3X�E!�3��$4}��2�����@��F��d�\�����]�J~�\ɐ�@�ɠ���x��S(/p�S��?R5��T7C{�y�T��v)�)B��tA�\A����k�ж���|����m0�8
y(��)����1UY��@�2�.��zށa��<�|l����\�e؊��U\=Ԣ"��a"s�(~�˩#������8�F�U��VUL�[I�_��ÒZ}��{_��L{#�F�~Ekn��Bd�Y5��Kc@��g�XlxV61EB     312     160@�����#�f�w��*�JB�Kzɚ�հE���4�����R	e����N�O��;32��6nRgj$��?�O�hPP�F��anm�3���_�CT�\�j(����w ��ܿ[7� sOk�Eɠn+�����#X��hA9��NV�y��id�J@'�OY:�0�%�E3U��^V����cb4�~bǼ�Q��0��UMj(N�ϑ�,�N��'g:�}L�(��mB�Lw�utI��*�LC*
�h�L�o���[���1�,�D��|4O�$���`������p����"���,����R���dTﻊ��-��V� �^zDsk�1�q�~G��:���^"'y13�