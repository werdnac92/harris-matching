XlxV61EB     400     130D9ɛ���l�k���G�b3�sq��$,�:�� ��n*ٖ�R*�Y^���8��S�C�ME���k�e��H�S�5Z�F7�n�0�nW�g='��@�vL�e�nm%����`�a�'n�E���h��T[�v��/U��#�߀�ǆ�^���e�=r�3�8�5�N3�2h�
?Sx�w,}�?�\�^����п}y�%8E�d��@��=�g���րO�+V�0����=��S���4�;�յU�o� x�'VЪ>nS�*A2�?�����fz����p�$eN?�+屈�ߔ�(WXlxV61EB     400     170&�$ǽ 0�Kt3���kFuÑBq���0%jY�D�IV���k�91 �eʚ=k����b�J��<}L�qDw����j���[:���}�g�������'A2U�`}����S��'x���Zg�(�)9��Q�3'�2����e��{��Vt��~�� �	 ����j��͋N�@mhDX_��h��2(u�a���:���!Ƒ�nn����;ܟ��ss@�2�gQd,�Û��h��!��#�{�W�5�t�����[c7^�l�oX`�!:ǽ�ah���$UA��������]w�W�/�'5�`y�D�9���=�����7�u1�ﵕB�d֧���Y+�����!��W�*��7~��q�����
�{XlxV61EB     400     120��0s�a�������>����{ލu��ҫ���*g�"����{Fo��.	�v5u��Pcf���2��f1}v	_�^��`����¼j�d�?H� ���(0�M���4}ԍ��X٤����o"�%��#������u[U��4�2Ӛ����K|�
^n4bu
0�qW�U�^��HZ����&�c�rܝp��Ujx��_�A2oQ�X��y�G[,/�0��@�l�W!hv��\���p�V��E������`�n���,-/�6߀z��XlxV61EB     400      e0�:�S��xiʴL/�V(Pʍ[7?�yP].g���D�H�I4d@&��>�A�u�Jڋ��H��<{��B���W�12��u�Hǉ�Ǐ�$�RZ;�0����?QE	���K#������v�7� �1��X6:z��ʣy���
S����K�Wm���	}�Y����vZ�86��2$�6�7��=�J�J�F2L����mP�������;e�-ϖq���XlxV61EB     400     160"��_�����̯�)�ʸ���@_�7��~�ߴe��P:��)�Vq�JJ�ufK4Cy�J�a�#�����s� 4��/�A{�4N�Ӄ%)?7�n���F\�#u���?�x���XV��v�U+p7�U�@2�2f��Jb�`���ʔ�}�����WDv��;�����Zz�N��{DI�p�G���Pǻ��1�K'�jקa>EQ\���A_��X�׹@w�s����'�s>iW=A���	e���y$,9�h8��;��Xc��s��c��l
����h(� �\?"!������"�T�&�����#v�&C��]�#۲�g�D4����1v_�>����/A��^u����0XlxV61EB     400     170�������n/߸��\\=��3p�����W�:^���%iq��kkr�Y�������o���*�1��S^Tp-B�!{��Q��,��������KB����Op.��^XϢ~�y1��)Ϸ�+���V8�x'�T=�ץ�w�·���DR�01�)����FO�^���`�n�/���s(�x^	jY/����$�s���o�n�ۏ�+���n��U��"���];���G!Cn���70L@��tK�o�A>��!���T)��V��Gm���hk������4�pb�4��C�O�rf��ϕZ���ɛRj�>�i�8�9!�vw�����1��]y��'���ze���>�b:O�8&��
�!./����qѨXlxV61EB     400     140(X��j��j�>:J,��K��I��~����C��e��S��@�2��*E����|�)�,��šh��:x����ʳ
l�ʴny<�C�
P��0���\�r�X�]��S����߃������|`�Ս�L�}\���\w��e�yL��������^s����]�����E���d���CgG\� T����n��*�T��(8-�w��d���2_��<����襁[�zL�γ��.Y��t5/B:A�: t��W�T90)#	�U�������Oќ,������t��
��`}�����@�E�[c�4�Q�n�XlxV61EB     400     110B��(<�������y,ho&\S8v�іb[��;���x[��ζ�g`7@����Ql�2|\�r_�"[��mp�݋a�nʉ��;�#x/��e+��׋F>��R,��>�lE����Q�ͻ�ohv���P�C5�eǿO��~]�7*��]��r��X�֜Gk2�l���g����9�s��v�2Ƙ>g�錓t�\&u�g�*�F¬i7W�Ks��o���J��R�O��a\\z!�����i���˷p� U-6"g(7�S]�PqXlxV61EB     400     130ĸ�X�����T���_�rU�pY���d�Di�����.Ih�b�p\� "����\Zz��C���u�u!���@Ȏ��o��E`�'v�~�Г	K����Y���^b���XCAK�լx�O����p�4��@[�~d$D\�ϰ���2�a�*�Ԭ�bJ�I�/;�0kv'g͢j�(��j�]�yĸ���勆��D�p:fh�N!�V�oV��m�.��g�XLQ�;����Kɠ�I�-������|�l$�J������4�p-o<�xYt
h�%�
��RW���n]�o ^XlxV61EB     400     170�A!�ձL&�o�m�
�b%�����'����q5W�1g�O�������[W�s|�.^ڱ�qo�����'�$�a���[ћ�O�[�W�N��C=?�[v�����,O7��N�M�\b $o����/U�2K��e��(��2�Ұ�m��h��Ft|��q�O�tN��.�#�mD�$��|mGb�J�!�l;����[� �^4B�5�P�lx�mg�'�Eg���V�UpFa�.�[�4F윤]���j�h|�e�e'�]8�EDb����μ��tt��S �-Y�/D)���-<������.Etk[\�}��|����ӥl�NY�Vt"���q����	�e Q8�ZɡS?���(ub\XlxV61EB      13      20�d��Dc˩�N���m��i]�]�@]m�z�l�