XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1503>���H3?���+iW��!8�9A����S/^�L���k�m���K�2nW1p���a��p��F�~[�?]WX�o��y�>���c��#}�FT�3d�����Ӹ�ge��3pU�S������d����gMxj��@7�k�"�m%���8�;?( %ۯ�%{[S ����[�H�H5��Ie���E��VGSEqS��(��&�1 ���J���Z6u�O�>�Ё��'��Æs
5p�ݹ�$(w8��f'~YϪ�J��*[t�&�~�鏢��+|�.�bE�J��y��]��X�jC��Ќ�<��7�+�0�4�3��.��ZΈ�XlxV61EB     400     110'G�[͋���_
���,ޕ�a��!�{+B�G����Ӗ%!fF�
�,c�G�����Xy��o�I�����ڿ|�R`�π���h���>�t�h�:��K-����J�W����=[	�D�+�N��\�˄;h�/�(����)��]�9�����d�%� ���k-PU,��,d�����//��H���7�kX�a����t#�D\c�Eh,�e@��W�7�n��_F�w��Ѕ���U�]�^�J#=���9\� s̐�?��b�Ǫl�P
�2XlxV61EB     400      f0�>��n�hao���(�jd*_��7^zja�X��n����C>����� 2Q� M�وB+��[��&y������2�����=!��{����c��nB��[a�e�b����{7
!:	f1�����A-kq�M��i�\*HL �ʕ;-��;��,���n�g�$�@�o�s���֢�@le�:߭�`*��!�tH�сQ`�u2]-�50G�`�~��=L���,��׀!�ļW�,<��XlxV61EB     400     130?�g[������v���w�V3���BOo~���L�ܿ3�+��1d1}'��L��8���h�d~|�g �{���*T�u�>m����v�&����,��,�w�
}�cS6)	+�fT��_����Ir��k>�ں���~��D!mF|VA�Nq�i�7�h��i6�7}>}�j%�z��NZTD�}��9��|��H��M�~���R��z���k"�h	��fX�9I_z�F��ķl<(y��>ְ�|�.�+#�s�2�W�]�~���6�u�������Y�`�!��3�":�� $=��m�co�
�y7�XlxV61EB      72      50E�91�s�`DJ�� 9�Ȭܿ�h��	U���HZ��Xv� r#����Z+݁��% t��,��"�Nt�J��U��Q~��