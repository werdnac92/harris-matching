XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     1a0�X�
���Z�v�i5S���H�|/��b����H���6gn�X�Q���z�T�I��6��IFn|_��n#�o�x���1��%S#�3'o$����j�o�(�l���i-c� �T˙AH���D�B�'�Vj� �z�~!�?���Px�'�\5�s�i7���tq�`��ywzMԋ�Lя�b���4%�b��ʳ�	��\G��oP�4{/\EOlی���+� g�ܑ.B/si�H��i[��X�c�D�F;|��B�(��'h��ItXt��Ϊ�-e��8�f%3��1���H֠���Z�Q2Y�qe�YAR�H�� ���a�y��px��\1 c�e5�'�F��iU����:+�8�l�3����ll��:p��V9�B�E�.}�t�r��RϏ%XlxV61EB     400     190�d�p�ܥg��vE	�UH����nE�ls:!K�2�`yMJDG����K�=�;co�?ǮX~{����"^�Mi�bZ���;C�I���w|�6	/�_4�űp��\��)s?6�ٍ���zq�s�	�Е\e�K�2�%��,��W��'ߵ1�/Q�7�v.����A���;���bE;ݷk�����\	���Ć.��NxfP!ϡ�؃$��xY���jk�c��Z������k�Ph����k��3NFɶ?��T����P��Y0W�~5�g�/�t��zE�����pZׯ�J��[T8���<�2E��sw���=Quw֏T� 9��A�Q���tVPTD7�N�A�Va�	/�g���FK����U�?9_���D��D�-�2��*�_�?XlxV61EB     133      a0 W�jG�?IK�������ߊ,�K|l�x����@,5A85=$��WAyH|PF�x9t��uy�,|1ˌ�Hv����vd����}C��P�Ks���nŦH~�@������� ҢJ2�Vq&��/^�q��B|C����2�J��:�̀�N
!E_�