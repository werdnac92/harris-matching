XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180-��բ��r�	�&w�Q$H�c�D8�:2a]��"
u�#$�r�ݞ�z�;\��C&���5�	Y���?�%����$EG��XJ;�e3S��U�}��K�F~��+=�t������ńe��W�,��JwM^g�coÿ�C�~����K���K��qp���$�c���+�:���(�EF:�DB��(�@���5�i*��{�,Iz��/pVV1�DRGl��G��CAU�|lJ�J�w�+�զcܼ#�P��|�Hql��J�H�}k	ho1�o0Fqe�W3>(���ǡ���^�ϰ��=�E�ts��4����d
�5��$!�g�ǻ1m[/c`��q���L����D�T�i`�(4+wG��'$A]�ݦ�ϊ�XlxV61EB     400      d0��/H�,����Pfn�?��1��X�Izπ�}����wԼ�Lu�t@�H]_��P��/9{0��q�}=�h�p�Sr�9�E���k�T20�K_��PY].�Ƿ�mgE�.����
��k狝S���$����kq�4��:�#�&E$���P��, (�:���:�'�h������u~݁Fv���؜G���p=�XlxV61EB     400     130��%,�U[X�c�T��38Y�	Q|���\ ƣ��5��2Mf̫� ;x�NKJs�P�63xt^�u�l
����e2�R�|�ϕ���L2�C�F�)ى֋���B	�P����1�9�idT�q��P�~"ݹV/�V�.�asUB^�A���m&��3��ڬι����f����G����	Ou�%*���0C�x�Y(r*�o������j}* ĬgR-5t��<K���=W���������^!Կ�F@�Y��]�������0ƌ09�K��8�m�mt��3�SҒ�N���x��3V;V�XlxV61EB     400      f0�n�2
��x��_������a�T���<�8K��M�*i��r]cM��Qeb��1s�
3 z>C�N���zߙD�Q�ё�]fϋϣG�3n�>_b �#?G����\���Ps�!5����p�z�I��K�GȷLy@�̫�!$j$�zL�9V�Y��+��R��tu?!��r�����3�@�U�g(;6�N�����ـ���.�P ���at�/�^Mkĳ��;�;lV	��ͩ�mXlxV61EB     400      f0���qyQR04C���N�:r�N��	�@���<=﹫��!�i��Y!fs��I���)�I �l�E	Fô�u|tI�%kO^{�:�I%<XA3r�#�.��O��z��1 �����C���w�M�]�l;���){=���i?AJg���A&+Sj�d o�_��!��f�J3��K:�¡�7cX������,�%���Lq:\�`HC)�ɡ'I�U���Ĕ�P\�n�XlxV61EB     400     130Y������	��F�N��$$�){&�iw�{Q�/�1ɟoX!�fyx���7��eNYf������#{ 5'���Műt�j��pV�W��/BJ4�/T�}��U!ϊ�?p
�clPoH�J��\U����т�J��b��G�3�\�i@�X�鸪w��\���ɬ����Zx>\ ���۷�La��k���\�<=,�An�#�^��$����4�A;)b"懥��]~�=r��&$S߈6�0k�s3*�_yx�tU)��j�*��X���<����G3>|�� uʓ�ٗoiXlxV61EB     400     150��(	2h��k���;T�zq� }�k�𸬺o���p'3xk����a�@�B�fY��J�K�k�ݗi(n_u/�wM�J T�#��!)K��}WR�m�V�h��I�˨=�X`
���h3g&�!��s�B��f)S&#$�l^���e��q6QO3���W \y��Ug
�J�!�}��`���=�&������-�*yl��'��+i-��k���Y?14��/���-LdKFsU�$��'�
X�)��l�l�S�����ޙa-ݩ�Hv43��ّX�T�_k���T�uyd��i�f�7A�667V�!�~����A����CaXlxV61EB     400     190ZO�����6��{�-�5��n�;��yW�N���L��^1S�\��)j��Z��sM%������.�J�7���l�)��_��</�Q�j	�ct�0ġ�-�S��] }B�W��߳���!h�����l�X��{K&EZt�����O�Ƚ1��(��	NfK����u�F�?��T�Dvͅ��d$h����	n��%�v�������3���Ԯd��A�Z¤���m�jakߨ���p	�����E�)]�l$yVs��tj��:��O�?�ɢ7���錎o\ ��u�ӒN%�4�\�l�H]㓈���d�)��[j�1�Z���Hd (�#��w�ݣ
n~���=|���g�@5Dq{���U[f,���׷�Uq5ͤ
&MH-XlxV61EB     386     150.�9�;{~���K�U�_p��A$�<���2�O"p[c��{�c!�;۠7M�k�-���c���ʂ��ϲ�K���ZP^���� ^���]����4�n��\��g�������.�'㻟��޼�-��׽�A��N��PC�{/׍�B=��9jcFoK����n.=8rІT�w0�#�;a����hy�^�6��Sh�~���.Y�LRjN��둑g �u$ei��q6��^Pw�G�0c�C���!���������:� ��4d#[��:�QFA4X\|��1�R�r�ri�����B�=�)��@�(��H��'.g���1��E