XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1c0���_�]%���멻�ٞ"q�΃@J�0_���a�������'�d}�x'zo�Gv"ڎ�sGc(�ۤ�f�׬K�P7��!�\�(��I���Ǵ�m��([�z2̺��,����R��Qw=�\X���/5����C���M��\��֔8�K���J��[�4���G����`"������F��:�~? �Bi6���`�>��ˣ��	�-$|`���������,�
oص��I��h�s��>[Z�\D������5�:l](v���ݎۀ�<�A'aw7 02nd�]��:���+�l5�� 4�Ћ��>��9�l���9���3���G�c{ʒ�e閌+�-S!C�0Ü[e�NLy\/؞�X��Kb�Yx����#ph�t���Ѱԫ}]�����O�з2x�=���PY����\������|XlxV61EB     400     170VQ���0��W��[u|�5IT}A]�A%B�j覶�eJlCb�I��ޙ�Q���-,d�2ŖsgZ!m����V��&��wk���J55U�~�0��ؙK��v��e� V��OA�+�r�1�a ���Ъ3l�{N����ׅvz��oO�n��:�{�Z��}&�7Պ#-��3�%jTdu)��	7 Y%�7?� @��
'�n�%�ԩ�Luh����,Z���=
�(�e���ٗ��#�]ʛ��aak���Յ�E�/�p�+#�BrBX9�S���p�fU#F���eu�O��P�j�w[Zhѱ�(�X����?�Gs���|��.����ߡv�v'o����^��ƲW���d��e�j�M�=y!XlxV61EB      95      60+�Ŧ� �qw'r��?�o���q�8	]@�U�[�O�!/�B�p�ȫZ# 5+�{��7u�l�:W�-�rR~���R��`�ۣ��e�Ç<�`�ٚ�