XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a0�Qc,�qȪ&�?����
��~]w�m!�΁�E�h��Y2?��a���T��3�\�!�'���h�dIE�)}�(f��2�+���^E~��:}��WTz��t�d4Ów�V�}�[���T�"��ޱ��ZI|�U� ,z�2�.�<��yt�S|��x��>��ϟ���l�B��3�h41	e�:k`p�m�ǺV�R���2�'���������T�Z'mT���÷�$�q�d��B�Ӝ�=dk��x+p�
 zz�c?����Z�<��v#7R2r��9�� ���}=@6X� �.M���}*�E���j������6����$KN�;u���\d��-��0��59r�4]���1�{�b�xӅ�(f��POi8��A1� �S�@�{�*W>�XlxV61EB     400     180���8P���U!��Lf�$�p�ڭD�#�U�-���5bBî:��m��na��>�	���7�R!zyy�X=��ۺ�^���*�W�b�uG�"�37v�����FFHƒ6'��;:џgÂ�f����r�V�m�Oc��yI�Jt�'j:B��]I-�� �}=��F�[_��iB�Czi�$�3	r(�K�pg�'V�:�K��a+;D�O�ypݏbj��g��ظ>m�0�+���'؊Ĳ��UI?��R�B9���S"a�G\�Ăk�P`��8M�`qq�\��nÊ�8~^��Rk� M�|r�a@#k�i=g3�*��2_��q�֥��ݛEI0��H8K箊�ެ���q��9�O6S�jןP>C2W�(KIXlxV61EB     400     110O=�UT��a��D@Z��찫��f)n�ȫ�lBX:v�]XFo������u�_��g���)�=y�Q�ƀ�g�r�{H�kGw��S ����_����-�0z�EX�m��7�k���tjc�.�+X{�� �oj"�k�;s�䦱d��H���__yV�eO@g:�a��w'�9�{E7C�a�l'��_��_
hM���`v��9t��$ϒ���`�� <��5]ֺ��&M5��b�����	#���a��1�ʨ÷�XlxV61EB     400     170,�d�b!Q\�0`a���a�;� ��s���4��H���/�Ɛ�H�,}��b���~C����qj��Y�q93-]{C�\�VB'�y�K�MzpA���5�S�W�ܜNB{�OS=M1�M�Ϻ揞9@ŔL#��l��ao"Q�0��0�x��A"�Ul
�ī������- ���!9�u0�"?f��p���>����v&.S?�
�q���`�llc�_#�V<:3�Ew-�,���!���gI����:.��s��@<Pu�29ٴ����,w��g]�<b�$9� 2�?g_U��Knr���=ҕ��I�|����F	:�T�_leBi�3k9�Ҥ�ŭք���[tG�z���%hϖw��OC.$�8.,XlxV61EB     400     140yM��&G��/�'���qT���������"��&7���߳���	�]ڌ����7�����Q��H�@�?���|���2c3�	�z4�'�[p����l!��:kB��㰶!^�Q�S#�<}��Bl��lѿ����ț�_�I�n ��`E���;�C��tw E"��V�EC���f�O��flęT��z]���	64�.��P�s�Ɖj�%f����IE	���>ԝׅ�;>j�����!%�4w��鞂t$�S)�ֿ�W��V�J�ʹU��#��%��)�s��\W�kH,~���'E�[͒f��>��. I��XlxV61EB     400     170U��_�H3�a�9Ѭ��F���#LЌ��^��$8����nfkN�6�]�G����r!l3�^�<��ד�U{η��j'�f���{C�ȿi�^7&�U� -�D��F�	"U/���:�㍨l��L����˼O%��l�:�0���}�&��f�:����K�wL��[��E�]�	�ZsS�}��i���pef�Y�^��I�s�.��ˁ`���v��G{�@أٟÖ˄Γ���6�4��}k�?�Û]�j�nW�`Hl��]:)��9=�^�<w�Ȼ��f���Ԥ�E���k�qq�l&N���!�xޡgQ��	;ۑ�#�J��"�Q�������o�jRP��7I��?lXlxV61EB     400     150���>s}a!�vЌ��VFȼ6�A.���������y�Uг��W�ق���aq_#�(��h/v�� \�)��Y�x�&!O����ŏ�i}��P_H"�<~��e#c�d�P��N&3�g6�a-+�t]�U�K�w[A�O����@ �ʏ\�%o�%�	[���ÞUF�<T�s ����9
�����Sz����Ҷ%���Ӡ�������6��}ӵp���81(����K|�m����в�z]��#6�锤|�4%W!_`��Ы0�3$�-�W������IYj���(��}����s�LU�3���'�M8jA�[	�W�I���PXlxV61EB     400     180[Cp$�����9t��D���U�{��%��;{�N�y��yI���r��-�n*7�!�3�7�V=GH�)׶�x��T�^�U"���"O�'%+b;"�ܧ�D�=hpˑ+��f懲���Y W8�jc�*Db�~^�������O��n/�$�X�|5����V�J�*��4s�6���Ϡ�W:!l�!I��:��q��\���g�w��޹��}���ųT5�M�����0�:�oX�XS�I�O�O-�n�A�ȗ.��j,u-����F������y�������}��4iBXe�c���t��(%��>[-/�<�4r�"hc�o>�Weñ�2�^���F�9�}̚�at��n*$��kY�P�1�W�XlxV61EB     400     160�#�kP��1M$r�饜���wHϯ���R:��9�|�R"pEW:�r�r�V@�D�޸���Jy�w������*�#H�ti�t���������!�|���s�l�b �Mʋ	V��8*6��f��Y՗�+�^JT�5�Y|T���EҚ���&wm*z�uX�au�����3�W�z���ێ��7�5i��W����g�ƪ����"]��)0���(`�1���,��w�mz�ڸ�����P�E��^LCO�T0<�Ap�U0I ey/���E�A�7##����]&��o��a���|�Z�U���s�;�Vd�g�.�І�ŔEJ��s/�dgT���r�V��z��nXlxV61EB     400     140�t�}���.r�=���$GD��%WB��u�`�5�_0է���T��	��nlJj���Ҝ^-t�	��?#A�tst��F�7r�k���2t�B���׷�F��x�\��f<Z�8�EN]�Ƽ�!
�	�=8�x6�+�� �ܜ%.N��[�ݔ~��c�|9m��!_�}H��߰�yR��z���s�k���;T$5����!Յ�z©6F�CB	>�h_.<�I�(O�|@��c<�0������w�UՌ�#�0�)T'�0.ȍ*:���RV��uS�Bh�Udk�������dSi�ZRF�b��s�0V�%�J��XlxV61EB     400     140���(���"6�U�G��`%hB*~>� _h����������g�{p����W��2�l{�ӥx��ws?�d���Y�oB���:���7�w��W*��}��F%���C&�W�����O�D˶��dft�*،�c�+�=�@U�p����R��_�OL����/�=�'�� �5i���*7�U[K������v1V&!�-��_����!j�z \g��<~����i�K����ֺ�^�}>�2.O6j��8A$}�S��X 0ͦ�ߒ��ی�yC5r6��O^�u����r��O  ��aA8��C`��L���q����kXlxV61EB     400     130kk�1��g��*����GΟF�1�,��jvH�ܙ'�j0�����(��I �n�:'Kf�%c,&Tl��IL�;���%:���#���2��@Β�O|�u��-v�@S(��}*<_����Fc⾵�"��V�l�]\�|VF.0�9��#�GϠ�W�
��׭[� ��o_P���<
���4�`Rb�:9=���X��=��	�K7�Պ�<zl�t��*p@��WN���d4�mOі���/������T-�T���I��E[NǕ�R=�C?i��>���z&Q�u��Z (��XlxV61EB       3      10Q�=���z�Le_�G