XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190��ږF)�L# ��G��i{���sƲ���k���3���0��ɝv��k+9YU��;���P<~����BR���a��E?ei���U����C\�����(�RU������"]���3=���W5��Ο��{��T��B*����6�z�]xY�}��{C�����q���s�*2��+l�,� ׍��[
�I����J�����y�Ҷz�~���OO�����1!˲W�Y��9����Q�{�Fp��� Y�Ɗ�zLb���$��r$tu�}<|В!���bYEP�"�+?`�s��P?���&Xq��I��5ݠM�3��ƶ���}�LgHki����G�^9�o�kă��2 S[��r�V
�DH�7s�ʧ��.�g��#�'��u��XlxV61EB     400     170�����Y�_S�Q��j:LK�B��AiZ�^\x�;�#-��t�90|�̨�bv���-�⫒R$�;�G�y������[XT=���
G">��ҍ�p5��|��;Ͱ �
��zu��:��)��0�tK����w�L9��4w��"���yx��[��Wu���e"�4�눲��q���5U1i�nO�/.ړpǴ�����I�R�yw%N�1�WwB�5��2�� ��6�c�J�38�X��'
�[@8/s�DzkƓ6�au��-�Bwȅ�C̖R���{�ޙ���$@�V&b���4�$�I�!�Ѣ��Dl~��, 1.*��E_��)|�,��6�)ܵ~$����s]����Ѧ ���XlxV61EB     138      c0:�?RZX�-�BY"�}�u:?D3�%����:�A�{��kK�m$���C�ܰ�51�t��\��b�UH����q��'
�0�u����]PBc	#��f7�
��Y+Eb��Pn87��fx���:!�ow]�y)�k�+���:k~}�SD�#ߎ���dXY]�S���8u�<�$
@���$��