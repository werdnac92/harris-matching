XlxV61EB     400     130���v�������b��q�`�������H�?-Gȶ�\�(��i$���*�����B(�J%��](����[/���> |,<���K4�2��4W���[ћ�x�G��n�l�<��Is��uGHJ܀W���nAs7�V�Ծ,��^����G�n��)�VR\�\�����AM���.�@�{i���o���������z����4O��[r�~�� %��Z���.Kx�)�:�y��h!�5Ӷ{���O8u�z�qf;�. ��5���B��������K���u +m�&�G�x%��XlxV61EB     400     190�v~�Y��Tl��;�c;�8Q�3V��D&bs.y�<��2��� *R>��[�|S���.eiP��r��e(�� �W�ɚB���P.�������v�	A$�+ǆ6�	��!�5p�pj��F�(t;��N�+VY�okE�]��)�-/�C��F�;�)L�hlʷ���^_ۉ �_֋͙��](YQ�NM�-|K�Ys�����G\iglОs��o�l�DܶE����r�_�,�X2W�y$��n���'�՟&���N3ƫNk�i�[Y�+���FlGTZ��sVޥl��M�/�؇����G��8�V�H�%s���	I!�+���W�`߃�}�����i
�s�H�Q\X��4�8�q5�٘�5N���E�B
��i�y�a��M�������!#���XlxV61EB     400      f0��~��hDM߃n@�s �c�%�8@�b�u|�e�������ځ��O�<+le�d�P��lq���0���	�q[:.����l���K��Ո�}"b�DF<=,O?��t��t]�(/Y/�nL��Cv9(�g���y㩕�bJ�7�e�~���^�X:X�Y�����΄A�8�᪙�EAP��4��
Z|���!�ߑ�6L�[1�����j37�'�xI��U4F? �j�A�	u��XlxV61EB     400      b06M���%�b�k�%6�yfg�ѐ��!��6l1����ID��@ei�7�㱹Y�4�6� !�{`C��q��<��~��]V���>Yr0���BX���t!(8���#�����~�x�4���n�A*��d���D��p:���'���x:�����rz����-S��XlxV61EB     400      b0_<&Pt��2�뺛:1J�O f����ׅ��4�O���%)�m�)㿻�;���!͋ٚp����6�բ��X�����4��lj;����MwS�-��a\䱚X'�fK�cFע�|G��ip�~�FUV;TEq3'�Q�1�G�aO8�Dg��|�|ᛒ
�V���`��>�����%3XlxV61EB     400      f0	�g��Dt��Y�����@�[�S�.\J��eF�vb�"J-���t����F���T�֖�Ѡ0��?��k�vS��g��.�Z�N쨉��&���X<)���TUs���w�R�ufH4�6�N�fd>��V�:�x����]J�J�	E��Wa����h��%^~�6��[lH����dLXy�0����Qh��DV�v�� Y�
��zYZЊ߱�S�z�b�@=�_�U%��0�z��XlxV61EB     400      f0^�ݳ��m3ˤK��O�����0v@	+>��S��m�&M�����yB�U��,u!�j�bE�A@�=X�� ���Q%֬x�X,h<�0 o9A;'�MV�lT�(w���M�rC��A�*+8��s��;�?�M�l�w���ɸ����S��Q��G��8�[�^�b� �����b����ozZUJ^� �N�?�0�k�Ҵ����:���+�rd��	���-,�X�g^*d�]�'*��?���XlxV61EB     400     160D��q}R3�c��,G&%��r�~�&�}��u�b��pw�u�T�̋h'��pc=�˅����g.�\�y����� e�"��a�	�	���!�$Dzw]�;�����r��y=_�.kRG�f �*-�ؤ~w�q-�
ݒ�YA���O_�M'y�}M^a��ǅ�G�S�X�3�����"�����EaEmh��$�8-[s�h���V��)oE�ߍ�ybH�)$$��=�s�SU�t��+�KeC���]a��3���z�W@�T�U�"3%��ڞrw��lRX7������y��7���a��U�/f�L�d4'�/BT��!<r�����ƪ�ţXlxV61EB     400     130�2�R��D�����x���Mϼ�"��eN��i���n�G���������QZ��n�.U�־���*b/t�p����g��uW�*�yb�Sr�#��V��c)ҋoH~ �J��&>#'t��G�͹����&��ǽN8�����2Ky�S�r�#{7%��E�O�˯C��ȜC����9�Q�w�Y�$'�ϬA�����៙m�q����d^�Լ2���F��y�@�
V�u�D��pH�f���S�"��/�E��������[ �&it����s��f���y!�B�aY�R�M�BXlxV61EB     400     130�.2[��zE�m��%l+�A��a5�Uf��(u���%��CA� {��ء�Iɤ�H�/a4��r�b|����vݨ�͎]_��	)�1z��X�D�2�s�#K9��Sɸ$��>�z��#�aOw ��^T��?Y���!1���ĦA���7��U������H�,7�A-�h�\3zY����<��7?H�7#��F��Hl)�B:��Y�^6�>���x1���gJ��6��|:��|D9�ӈ���ic��z�<Ǽ��i[��=9��]�:�{��è���L�6��D>v��<���
.��XlxV61EB      74      60R��z�RxRG&���MD�u,�пG̦����9뽴%�If��V���
��S���Pe�v����&~�����4��y���bt�~-vAA��Z"