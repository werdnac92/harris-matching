XlxV61EB     400     130?4�ی�X1- uǨ�
E�>��Q:�H��Y*`r^>t���t�:�㑰O�%��w���M��%UO=��1T�?(nl�x�|�qY�>-��g�)2oN����7P9KF��߁��Q�[���i�����i�qNG�ǡ{"J��3c��M��sD��ϰ+T1�
b�y�˲0�:�:=��i�	�?^�nP�'�����#ޥT[�ՃnD���j"t�d����w��H���s�o���~t��os�<�w�������<��튑�RrT�x�M�y�Q8�
���!{)
��+l�W�A��XlxV61EB     400     1b0�D��ю�8�m4�.�j(�
 h���?�we9���j�TE�[g�7GtCه�z�h���h!<���w����t��N��Ao�k�<]�-��
�;�"m����Å��A;Ob�>��������A�)�)-�'�A��P��u�Gg�!n=�"�$%�sTV����z����r�����[�G�!١b #�o���l��w�L��H��5y�|>_ �0��%�����US6�uH��N8y��?��)��^���\�+		S�l�pC	����/::���RL	���YT6ğ��^�����L�)����36���~Ja+�\i�W6 jt�,]y\�bvg�j(�p��@�����
����@�AY�����{5�7����oK���q�Ƚ��Xh7nW>�lNć����Q���>S[�XlxV61EB      c9      80.�R*�3Ԗ<��r�^����?������s5��,/����%��͎ɽA�tqq��>%M�:FxK߭Е�6�ٙ�����O�*��Zw#][EUV��U��	�2�7Y>�n`eñվ�$��