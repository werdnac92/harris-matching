XlxV61EB     400     140?4�ی�X1- uǨ�
E�>��Q:�H��Y*`r=%nE���p��b��g��~GudST��)D/_�ߪG1���v7
��О�l�(��a��NUƿ��a��D�����]�(�=0��}X�?RU#�
rO���+`3���T7d$;")N��^��O��㣅�����[ظ�{WtSK���-t��pD*5W��˷)�rs��v�y�����Z"XV2�}�v�\ۃ��<�T�n���� Q�� ~�$J=�v4��u�}/�A���qCt"�^h_vO|��ԩ��i�!=񎶽����V|◱����XlxV61EB     3ef     190���%�sw����@�$3{O����z�)��a#���kB)�����y��È�����MsǞt��2�G�k���)��_��I+e�nV#xw2%��\�<�Ij�+͊/x���kT/'��OQ� ߾�i5��O֤�d�D�	�I-�����bc�;�E�o��!<���Fd�D���!��N$�R;�v�z7�/��2���$8|�g$�@���Jq����-O����b��q��?�-�b�}�g�N?��4��T�`���L����m�9��{��{?j�j���E����vS���ɱ�y	�Y�:fc��m��NJ)>�4+o�	���J-�Da�&~�ɡݱ�w�4U^ۏ]-s�#���%U����ǮJ��I;��c�5c0|+�O�8�ד