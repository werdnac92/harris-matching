XlxV61EB     400     130���v�������b��3�%>t�*N��mc�r-���>Se�{[��� ����p�,1�R]���;�gxX�(�٦���K&X��m�x��4�3PX\�b4��aYn?��pg���jYuj����i�
������n���鏡D�6ե���S�T�����/�8d���Alzie� }�ʽM��&���u��a��^meL'���Hm�I�yV$ɀ�ћtl�s�x�b�@�eX���|\A�[���[(���2�Z@[�f���ӝ�W��Uh�!�C�E��Q�jnd-��{Zv�XlxV61EB     400     190*`��FX�	O4p��� �s�j�9w�<yV��������̄	�Q䬉���a�g�v0J�f�:OF��i%�$o3��50��t���^�D�E��k��̀ڙြ�b�{�]AA8MG�:�2z-���x8��z����*h�����6�6�o��:A�5�~�hp����K)`$isV���ô���q�|w��ƭ�}?�P2ow��iŎ��-��(��e�_ǌ%��|K|��~~<��i݈1� ��f�I1*%���Q~��^r¹���ZLb�'��˩��ˈ5���]�4�$�ȶ��[�ی�L��5�^���i�9�?��1�� �w�A��:J�V�P�3���{>}0��"��n^6���Ɛ�c<$+�aa�=9���bXlxV61EB      c7      80�^u�9��=q�������K�k�v��n^��&߀Y{�RPJ�%o������2F����ѿ�&��$��ٱ�V�׷�|W��N�����|)�:tp���+�i��{����asxK�C�q7�E