XlxV61EB     400     130���v�������b��䥰-j�lM�K&UR���~-�܃�M�۫��F*�ɱD�@��>;�y��*n.^7�'�'��S5��"�����u�����FYJ2h��yE��;-G��.��+-=Fm���{���@��!E6w
{���G�y�=�A"s���"qҰP-��*s	����;�7���݅f�Ś�c���5=�çi�A�A�T���twaf_�W�ME6�K��2h�d�L�(���;Op�0�"���u��,. ��t
��W��uP�
�Յ���Q%��(W��@*�b�s�+BXlxV61EB     400     150C�m�P �5�w[6����bG��CX�14��/j�%Gw2pQ�{���44�����P6� :�6��6��f�],2�3	�M�\��aϕ��ɑA�v�C� �92O$�p��ϚN��%���(%DӰ �c���e遘�U�G|�
D�&;��470d����|����o��c���l�1A�0�I���a�9PW�c���R��D�X��������]�q�u:ڱ�(�< .ie�n��'��X��s��> j®U�g��Z�c%�N9��2��D8�J��#_��r�}׆��:ݢ��l�-cN3x�׎Q�.����"�	{^5�6,o�4XlxV61EB     400     170��*٠�k�28���$<����6��G�P���?�����z����\��b�*��}��rк� hT�&3r��X�#l�Z�����0�_4��:>ă*���=�(@)��rb�3�9R��P��_�`�(Af�A���va)T��2��)�0?yo�G��g5�މ��a��������[�l����-�7q�Ȅ�#�ض܁�cT/�����V�)6�*����w�)7E&z�wVEH�������eæS������lڮnL�DJ�_*�^�s�~���Q�itE��ӞC\�k����9T���pShA�y9�ܵj��a�2�#������&���yHƓ���pB/{��c�<}�C}�{a�F��L�YO�yXlxV61EB     400     170k}n�-�e�fSJ�n����y�\�@A�6,0��_<��
7�	3����u�f�����C7��W�v[u>�\�n�7.�/���*=�h8��Bb�s��T��m1��m���-�X��w�'Y�T%_�ž�qPX��ƾ0�+�d7o��*6��;�J��o	i�{2ir�
�)�h���|��ށ��M񩈓'�o$Y��;ٞo����<�m#�)��L��>�WAX����&�"�4A�QJ�[�v�':����}S!�d����@�6�ϥ��j�ŗ �u�ا���U麯A%	�:��`���>5�A�� �!ׂ��E7pL��=�x���J�J�BJ��.��I�K�GXlxV61EB     400     1b0���1��/��%W����L�;�������x�8v�㭦��!�	{�����ì
c�K,J�~J[��3AKm�&�FO�%���DZ"b'��>+<޹���_8l���5�.���j �&�ױ�mxn��t��v�6�h\'������,��
��4psG�[b��
Rع���+�.�B�
����Zd�K��`�T_f��e��}���ح��r����� �0$�9:A����� ����\J+�|%�q���U}n��R/XXYe��Ԏ2�VQ<<�.��ڂg��W$(�UXe���U�IN�|ɴ�[ك��(�%�/�3�5��FT�̰�ʉ���5E�U`;T��m�&i������gXs��s�X��w3C;W461i`}X�4��9M�:������͊�����:D�:�w�Y�<������.��+�XlxV61EB     296     130��!�� ��-�x.O�T��h\LƗ	7�٥b�����^��7?���A��6���l����2ٜb�T\�v�;�j�.�B>�u!f���f&�u���m�^��P�}Y�:�S�<"+'��mٜ��bMd�	�ħ�*��By���u0T�m�D�S�b�����^+�Q��M�������e��
��W�؛���;��i��	�U���둔�������&���&?�Ak2�Sdl}!�ܬ\�� �'#>����}��@�g����9Q�f�A��q�8�]�OlN��v4_�<�