XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180P�@'��Z���]��N�	�K���\�m��q��zA��ゾ)�ێ�ev-aL�])֥�w���������"�k|̛G���|�{���+�46�>�׉P�i#l��V2�YQ�F�J�R���������Mt�~1�^0��!6h��p��z�3��H�'x���pni�95��|��U�&��cI�񶦣r,��ܙ�ƈ`D�/ˊF2q��Z��蠟�w�=�����u�
�u���Z֡d鷦�<#;x�^�O�;��嗦ơơ@��lZ�������ѩ9v�#��K�`mxLV.Vp֩�Ԩ����K���x-��Or�8��� Y�qv�::�7	�3�U�kIWB��rU)[֕Q���ּ�$����=��KP$�E�S$���XlxV61EB     400     1a0��.���J�����Q����ۺ���ttJ�M�.�����A�F*_�,�Ǐ�y|��H�#\t�uy
��_��y��U��oF6�c�a�.���?�Sz{�\�-{^*�qLv��fT��Q<�΁�*Xӏ��0q��N�>N�JU�2j�$;�z�j���0�0��E���V���ׁ�p)#�?���	�HG��2��"�j{8�k���N;AUQJ��l5���} �#Co����.VG4$W���-�8�lǑY������lc�w�B��%\�d C�GgH�
���օj���ꅸ��[8�B�����p�Am'����Fѫ�f�2궁��>u ���I��븴���̳�ׂ�w�y�����Ur��1�|��[�� ��׊�$�~���$5�Z���m�QXlxV61EB     400     140TI'���#���л��Cɥ/P`��g��㤪s@��K9�F��GZ���Cg��|������Or6U��0؎#6D���.�(��d����P�Fۓ�ݮ
p�*���f���i<~�������,��Q?��N���'($;d���f�c�\2\s��ͅ0�9���,������6��J�V"�O{\�uX\�mr��?�Y�N�l$���1�����$�>@�0o�mmCEy�[��g^�<����q�\��'�hf�	h��p� �����u����X�6�={]D.��k�� 	�ן�H�	0�d[XlxV61EB     400     160�!T�C���G��ċ�&t/L�+X��4R�?�kҍt���B{��o ����(�u�^+�#υ�� �,�|�����Q��)'Y^i,����I�<�I�A2}�{A�G����/�	j��G�	R^r��$I7����̳��9yG��d^o%ڤ�d����޸?�:Y�"�B��� ^�dws8�޹b;A\.	LF0����'�n��D��G6�@$G]5�օ]�)G�l��ۂ�V�A��0Y!-Gth���A�^�-�I�v�jy�/o��	)юW2��L�<��+���1LBK&`���g��ξ"9АosE�}�>Ѣq"w��K�2��d�+���RԱ�T�+qXlxV61EB     400     1a09��rb&Ǳ��t}ˈ_C�����b,���s#E$�+M�bn��Qs�B#�U�2p��� ��"KG�>�m��X6������k��T��X�ڌbc�|1��K��a�}�/���lx�Īj��}i(��x�R n?��D�5������m�%7o$�<m�C�g_��-�n���/*�t���f�du��Xd�c8��U�**��Hp�>�������8�MI�8��5Y��˅f�,�q~y4�9w0z�����۠��tJŌ���.���4�*'�+����D���y�K'���	[�V����R$�F��><��7�r���֬�YN�.
]V�-�( �1��[2A�ZA��B��D�?��ʁ(� �g��:��vQ~�<�DF��$���{�6����XlxV61EB     400     180"��M�LH]�|f����y�������[��Y���O��N`_�/�5�ލbG��	����	��1a�=�J��%Feec�[hQ<P6�H':�N@0�g�΃��W�Lz=�|����m)<��;�o�W3V��%��7��"���+
�t����B�g�]A�6*6�n��ݺ���[�[���#d�e�גr�B�+bLh�f͜v�)z28⩕.9�&N�����ߴvX�To:�FLn��w�\!�bGr�y_��2�0^4�02���l�h�6b%'W�+�K����瑛�U����\W��Þ��"�x{~�+�_XYP�g��C��R����΀�r6�7>��.ݓ(1�&��G���hM4��K����XlxV61EB     270      f0�?��R�8�kA}�%�.A��������
�:K���L��~�����o���M'���6vC����˺����~��U$��>��6����vcE߀F���>'E4`1H�ݒO��Yܳ�hi9� vw㴲N�P��xb�*�A��aB0~����/,�_Q��R�	YźJv� }Mjtw�黗9 �jM�H�V��ʩ�x�����iI_<�9����c�R�3���I|'�Ư	D6Q��6