XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     170��Y��K_͝G�r9��cxRM*�+�)�IJ!���j����x���NA$B`�A�Y�Q;M�"kJ�f7���i�gd�6�m�ȃ�6;t��pJz�����V3���.��T��d�b�z��-�� W4�P�������Y>M5�	t�^v��Y��)�k������sĿ�d������=��hX��-w���ҫ�a����P{=���}O�����æFy���&����H��:t_��=�*eE5|�]�1�3)���m��n��̣r������`�w*����ul�����x	��Ć���t���	���;�!%)�qDI��<ݒ�{����M���q���8?�����KV���(j��f<i���mXlxV61EB     400      c0�+���8�QP,'
J���UR�ӡ�|l�X�Z�Ѯ$d��_�F4[�5Lk�.�Y��U7�#�����6<Z�l#�c ܆$�pl�� �OV��C��3��NZ!��;0��,�)⩍Dfh.s����<+��%��ౄ���
��?���D�&�_-`��	i�F&��5R1p��099hXlxV61EB     400      d0Ȭ�Qu���1Ĉ�s�Ȫ0k����76����=5}�t�9E����ޡ|+���[]@j"3��a&��"�0͔���#�K�� �k?Æs
�)5ԀV�ˑ=@�ю'?�d�s�#�\���;˃/+a��I�!6�u�'�dB`��D^�<�	�x���"�sᶠV)|�$h{�+��t���n�U����5dp�ܜ(��<�ʁ>Y��XlxV61EB     400      90�<Y��6���D��AD7u�Y���d��ؚٻߔ�d��%�ǂzH7�f(u���Y q/��g�~��\�⥽����M�:���%΢1E7�YG�IK\�����n����y���;�>��\�3�����>u�}XlxV61EB     400      b0FNmQ ��"6���@�G�os.��,�8�g����	���,�Xy�F���v/d�w�+���9�{o#���Z�0��,��0&������ ���Ja�&b�"��)�����ݭ!��g��[5��#��H�8��x��X2�(�S�}��z1e�{o�� �:�aC����:�rA�XlxV61EB     400      90^���ab��R�d�U��M�|EY��D�܂�<��g�'|�&��0� �+�� |V�q�r��ߪ���}�J9�����Xc�:���R�ba�x�#����l�[��_[��x��^��s#�AB7���q�����Ay�H�F����o��XlxV61EB     400      a0���J���P��{Qܯ������Ә�ʧ)H�O<1�x4W����sG�2��L��&��� t�z� (hz�kPYL��L�����O�'v�ʚ��_������t��Jlmf�o�7����M��y��|����5l�v���|��B��"�E��0>��XlxV61EB     400     110+������l��ӽ!�s��RL����| ���p
�����'s�'�=���d���\l�f8�����_�Z��4Z�@�� L}�'��RH�ɬϫ�fGK��+([���.J�m�/1$[k�T,K����q���brW������)���0�vB�a��b?�b$��dRtR�uO�Li�l���	��!��"^�~���������FH5ZpN��5on���)�.�M�eR������>��!��������T�G:9�Um�� �滞��Hg�0��,���XlxV61EB     400      e04zN����՞㯄�\~M��Y13�[Ec�gcvi�����zNSA
5�50�T�6�-7oed}j���Pգ�C��Z;�y�)���NgG$ˀq���<��x���C ���+bZ»(1bn��v�ò�ϕ5;�����d�T�Kjh�[�	~z#�,w#��D>�eݐJ���51�tՌ�v[��"W���$!��V��@jT~:��O^S�Ry�&��`W�4�P�XlxV61EB     400      f0�I�k�;q�PXh�N��*%k�����{��X�` �v*x�Pן��@��\K>�3[)ߗ_� ��
o���t����K������_��F<�� �}�oN@Tڇ
��|@�!��vO?sf��z i��O�r;�D�ќ��<ҳFH���Lhc���dC[l�/-��h��^s�m���@��-
����D�!����~(݀�d��L���:��TN�ʋ�B��#�~�0�u�&����w*O�XlxV61EB     400      e0`���V�4��?4�deQ��/V���4�-��
@��/
���+�H�p�1��Hu�a(�TkG����`:ee+v�"�j*��xX�5�p�	���0�P�a�E�aL��D�:*L��6adaٟ�����!��CH�����r�y������p?èK�� p��ڎs�4�����@�=��D�b$�7�v���VԹM#�G[��<�K	8�:�P�-�	�?%�ΚXlxV61EB     400      e0x���0��j�3?
šW�x������U��6�%��F7���Z|ϔ0h�O:�-���i:&+m%�GF6�Z3n�/�`��q�`��������������g;[�=�t��#~N�1�;	�Ƥ�"Y)R�� �|����\Gխ��vZ�?i=��4ƽ���S)���E��UA�/\(j/Ze���Pf�����P� �X��َ�GJm[܂�+U�4 �bD�`XlxV61EB     400      e0Q?!�9��`�Hl���@x�աU_l� �"m(�l?Ϟ��ʑA/ٮ :E��
���)��~�<�޵��Nl��ai����t[�e��d<�����궛�Qz�?����-6MѺv%+4�K�[���Y���0�����e�A溘5q��)��L���-�%�����U��p��7�3}s[@Qf�	g��*W�=�s��j��[���N[p~�c�j���>�q褟XlxV61EB     400      e0G�awn�'���.fEr��JAL�'}p�$� $�'�K#�;1�[�A�پ�o4�:ˇpȉ�� u$ ��/�ǵ��S���&�;�X([�HҸ��a��w�~GjqI�����ec�/�Ā��=g���'�������/#�;�P:�V����;�x��y�tDq^	-���Q�5џ�_9t�ӄ��ş�l��-|bA��M\�jNz�\�ޝ�ꨏrAXlxV61EB     400      e0HnQ���{6b����]�C��^K�}�x��8D�+�+�K���L���z�d.�3>,�tW8x"�y
C�2�A;�AF|x|p��A���*�o�vg�fѓ-A;�C����_NQ�O�2�܁;�G�qΉߤ~�v�^v>�.��K8N��U�~ΐ6)ɔ�����ϒ�78>�$q�r�R��.__�(���FQ.NR�����zl`�Ҥl���~��XlxV61EB     400      d0
�VX��pU')0�;2�VW3�?A�]?;2s��������.�`��9�r���0������AX���z�c�q�	v�j��\�c�EV�#?'9H��؀xZ���]�&�"��Հ�m���1 �\�,��ӧ�o'��}�LC�̰+���7`'2��0�=��t�S��l5fz8K����E�,�fP��.u/��v��t�Db�&iXlxV61EB     400     130�:F�����j�y��k���)�m.��Q�〔ӏ���{�,�
��`-=��m*'���	\���H�PQk�m욈�h0'�sd�F��e9~���&Uθ ��~� �"����k��J%t�k��*H�]ɍ�hm����R�V@��P(�V��(��7�JպU��|�f�����-�A����j���Ɓuv=�"�יآ�W楉�U[�oϤa�d� ӡ��{+��頨�����3�~�Hž�9o�z,���%�iz�I}�����|u��˔<MY�;3yN�gUJ���>8kXlxV61EB     400     130m��!KN5I��bT���y\u����{���rxnϗ���z�i�z��"'���s��P�����b�fϴ���m�<�ox2ۭ��	-��|<(w�v��S�e��J�$��`������ɜ����?K� u�� N���Ƙ1 �����C�U��Kd��8�̰ I�s�"<�$��^��)�,qH�KG��u��ρ�Jn,H]���0��RF�R#��� e��#�*�sc��~�K1oh�\�}���J��� �Z��ٚ8OU�� � ���xP�BߧH���<XlxV61EB     400     150
��W(UH�xO���P`��0j�-�iz��S*}z�1>L�����w�ܳ6�$:ZX�Vv'+�vL��mn%f��Vn�Ë�Ot��ϩiK�̤��G���*5S66��V�6����W�O���X������K~�.��M�;�	���W����p�ǉUd/�_�*�tAK� C�$?�)oE�������:�G�'�*� �
M�oXe/e��H�6�N�L=�e��g�+�@�7q`O�҉�o�.�L�b�Ѐ�#.��n.@Q�`�`g�dX�+Y�se����-\��x�II����Խ&�U��q�l�@���\� �@�����P㡛ѱ]3XlxV61EB     400      e0���a )�5�7�/�_�^y~+ˮ�b�5���zw�Td����!�>'%��bɷ�R������H�s%3pkmhL��e3A0�������r{:�3��ۀ�\V�����ʉ�~?��6(�� )����>ن��便����t$ �ؽ4@�L9K5�˷���0�p�xt�^}�l��B6����������m����)�d�o�X�w���Q����G�@�� km�Y��XlxV61EB     400      f09^|.�!�)��뛀�j�SS!�^������Q8��g%f�����'y��#���-�X� ��i�I�X�W54����j�0��(�� �8idJ$�@���^�
��E�g�KKʺ�#��b'��������!�#*�G:�������;7�w�9��=h����%�Y����g��>0��X�?��u�u-�;TiY����F����R�3*� &� /�ƴ�h�.�i�'�XlxV61EB     400     100��N�;M���C9�=4�^�
���5�M��P�����"�I�}eh+ ��{��l��x�|#�S^�Y_T{̶��{���{�T���J\T�`��|��ll�u��˅'�z���\��)'���)f��[F2���rKy@дIw+_I�@�u��1��XPuN�s��<ѐvׁ��ߴ�\A��]#f�����H��&&��x�ߐ���:;�Ԡ������h�pu-��`=|�� ��R4Ɲ�k@�}��@z#\�jakXlxV61EB     400      c0�
����YmCbMu^YӔ0Z|��V��d���~"L�n�~Y�E�#@���w�.�h�"A:\b��jdƧJ��ڝ��n�U9��=r .�K���;��0רn��&����2�[4N�d_S��2d�W��ZŻ?��b|�
sy�����(��ř�K�щ��C���yq�8��JRe��_����G_���XlxV61EB     400      c0�.E���sB�l��d=0�R����JTc'!�?��MP����o���+�I�qכo���M:I���,s������M�R�I^&�#wF������	P��`�Z��(Ł<�B�e�0�ec�6?����Ut^P�;�#�{�������_i������s U'����r�O�{|�c��ܬ�q	��WXlxV61EB     16e      90J~L���<,�o�B�E�Ԯ�������Sj�(}�hcK�/d��s�&�b�0i��FƊ��H���n�i���;��=j��9$����_���=)�)݋�������Pgs����`� ��gN�|�h<z���%�)��