XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     160]���J��� YĚ�R��v{w`�{?a���qɏ�����8MJN�w�Q���8{�}r�,���`j9�JZeI��r��I�_J-.������//L�wy��������gi�a!�|7����(Q��h��_���K>�qbZh�����򤬩1]�}��{>U	��]{D����J�q����`�G��.�U[��dn��P�t���A �z3�̻-?�1m-����J�ޏ�ā7��V���]�G6C���S4H���N�W��4S��.��F�1[؀s4��ιt��r�j'^t��i#��S7OQ��W裴 ���@�����:�<!XlxV61EB     400     170�`�݄���T���l�8���}ߨ�16����ƾ;�"��HPH������p�Fb9�TzD�,���91Cz%�Tr���t��du�[��H��	?���[�!G�̘�;���/��5���׀�d��~ʱ� t;��f8�!-�wr����tOO��Ό���7p'|<(��D ��@��l��y���ǳ��X��i��,�_L �jC�V�d��ㅋX��������h���\FJ���������I<s�Zwc�3��T��iG�~��<��<MXsU0�q�A��S��τ�]n��8I.C���m���C#]��=p�o.�w�v�X���JO���X)A4׆x�N�c(F�XlxV61EB     24b      e0p�C'���(Pr�f�����vdQ������%n�7��!|��&W�H\B�@]AFڒ��t�i�F�e�%��u|Χ�A�61���W��r�P9'�|=گ�Nm7#�4V���ԯ[����PVc��������q���U}��AD��_��AX��{	��������[	��ԍ��	��,�=��F�>�0��������uk������mp䎻+FG