XlxV61EB     400     140A�?7��'͆1H`�
T��g���	v;vy�8�D������*H��Qw�����G�������(C���x)�#���<�Su�0>��:�����!���g���elB��w~�K����o� <0�J8����@*��+_�}H\�ZbF9J=@���P_D����$O&6�����L�U;����%l�4�ĩ7^��p�L!�-3Wxpy���)�J,��qM@��\#����I�rx}k��Q��.N�Xw��Sv*$Vd�]��T��20���a��<�� �߃	F`�
,,"Z;Moy�e�5������9XlxV61EB     400     190�y�L��cW���R,iU
��bZ�-z:nD��>H;Prl��{ A{�����Ѓ�Dz��<�74��i`yGf�`�zZZ~G[�{+)9-ԠT3�����Kp�D����Y^��f��β�녪�	��e%q�#C����
�0tG���s�mܬ���U�������� ��7�`�$� �)۔v��]�*�M�5ٍ���r3_@>�^��f=�w���x��Ô�b��诗^���#M���!���f�h������e�WP���!��l>�ۿw�%̯�`��ci��~�#X��S�/�5��-�<��&Z��\�s�#�?}	�q��5Xacs����j/ĉ�'�g]k��(� �_R��\�n��\�U�����"@�N���XlxV61EB     400     180�i��P�?����p�P��6��WlT�0��1O�^pKJdy�*B��2+�r�1E�tT7u���rw���A��1F5��k�@�F�w��Qv����+�5�1�TH.�H��b�R�6�F���>�>?������~d�ղ:M�5+S~�6m��X�һ�2�O�]KB-��w!�T��Z����ћ�*�_�Ù�t=�P�����]׉�V�V�t/�ʛp�.	Y�/E�����eٌ!�	����c� 04��[7���>�j�!���2x��:�/A��c�▯(D�n�,	�)�����e��L2�_ ,�8j����De�r�w��6����v�sV�oجI�^2<����n�@���m���[�"�*��1�RMN�>���M��XlxV61EB     140      a0�F�@0�����/Ka\T9Mb���ʝ0��7Ʒ�,�;Fte��Pڐ�����g:^%TJ*N"��g�Nx�;�à���f&Ӷ�Q��Z��`���'[��"D��/kI��= $��b7���X��Ѫ ��a�>�fl+�_�u�r�Sx�[y��