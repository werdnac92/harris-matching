XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     160|�2�yNF�+;�(�PX%#�d��Ę~dym7�[=^��2��i�����U��&Y�yRc�T�!�i�d<�ߏ�8)��&Q�a���3]���k-���a�yo��� 7�+�	0v.��Dq>7������� f	3�0=�g�t�_��n�_� Ȳ�{���^�Ym���t\	=�+8�����a�OS�皷�j��$S(�^h�<#�rbkIR吷�f�[;5�H�u���$���;$U�*	ey��ȟ�$���N�6�d���s�ΪB�A��}�� +/6sEy~�����xb3�%-��>�M�=/'b��5����)��m��o�wR���F�@!��;C�WXlxV61EB     400     100R�k?�g�I����0�7m�tΓgm�?A��ff3GhYp�.:��P�[ԫ�i���]x���WݚgX�Er�O��aɺ((��?�|[V�\�!b54B�Qp�;]�]�|���o��j�3O*2J�ǚ#R:�ȥ�gO����j����D���:��@!��W���]N�B6�Dd?`�g��L�9�޳U�v�O�j���~!��r:���L�IRQ�5�X��wR�*W�Е�GvN���e��+�w�ꢣ�XlxV61EB     400     1c0>Ve��3ЉƄ������#�G͹�_{���zi4*����Q���-�(F� ���7��P�n���c���MrP��s���C����zULck�U���;e�M��S=�Rω>^�R��Et�ϕ�_+Vx�^I���eD��ȑ�2p��X���A��Q���_3�R�q˥�Sb�mC�"�:+9-����Vۻ)0�V��|@E���{ �>������Z��Y��*��ר�b˧Ugk��&%��'m�P�Q̟8��>�n�"�$)�<710�1��#��'���01�
8���T�GRGĴ۽��jv�����0[/�Ȁ�^v4*�tq�����+ǅ�uR�,{&⪈S�ܭrI�M�H){m�*+ D�DH^8���R)�����^�vI��/5���3�Z�R�,I�W�ˉ����3n�E�n����2�c/����{��XlxV61EB     400     180�/��(2��B���5!}�`N�7:���}�/�I���d-a�/m��hX��r��m�b��p^�����[Մ�Ɯ�n�v�!����V���/vgFK��,=!�^�7�#��'W�;er�����@�W3�Lz����������h�����:4����N��I�o��P��S]��J�t1u�<�����п>�gO=����U��s����<ח���ؤ���������a�<�N�@��G	4g��e����Ew9u0��z��Н2���k�3�ο��R�ɖM�v��j� ��fڮ��׏Cܮ������h(�6���( �5�
ôC
䥽�A#�42�\��M�,����Yĥ��lX�n.�FA[XlxV61EB     400     150�o�X��/��v�,�+�|ʕ+d��ᒟ�Z������G�a�)�+*��}�"�Ԃ�i#��ߛA �I���X�/�G����a�dNK'�� �33�\���a	�_z!�(��<9>��ޔ�6miW�O0�#�7Z���-آ,R���v�*�
j�|�Fs��t�>������$�I�����ߋ"Ye�gf7y����w5����c����'�%b�i#��7�F��M>?���×?�Ĩ������ aR
A��0��y��#���p���$X�R���vuD�}l_��N��d��4S 6:CJN��7��1Z�ՈTtz�� o���׺��!XlxV61EB     400     160Ρ��J�^T�}\x���bO?����������u���F���@�?���I�_�\圯��Z�q��_��~�Om��k�뜂�	���A�J�T(�G`RJ����>>,�L+>�U2�EB���=t�_��K2<�=x�'���7�Ԟ8��>�Ԙr�kr͸F�̶���w,'��ŵ"#�H�J%�ٸ��hi����⪺ާp�t�F����V��0�?� c�]%���0��b�hx�`�{'ʏ�-��L�v~�T38�]�_WC�9<��<�RU�	UEF�n ۃ��,_�<ag�+P^3л��0�ד=Z�<�,{4ΖU���$�]3j¢�h/OP��$�P	�XlxV61EB      31      30V-�W>��)2=�z_5�44"���f�)W��_f��elz�FO��