XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a0�?MϹ�\�J��=���}b�-i#14	y3�X��V3����>�N��+���zO�z�@����E����j�&�VE���<M;g[�e��7�	G1쒛'}��w�
���2�l��g���M#�o����h�����U�ME�8Ͼ�P$�7�z�1X�m��{Y\�o��?�5�o�Z/ �1,d-0G�9U�9�����-��#�(�79)	�JkJ�g����ٟ�hM�?ݷ� �L�T/�Y3����յzy��tm���7�C��@	�G����� �-gW��r�}K�_�CUj�8Ӗ���7�=����H�,�˞D��^5z4��Q�qr*]k���f�n�e�=��.�R`N�щs[8T���4��! uM�Μ���j����e�RO�ΤI���l�B\^���XlxV61EB     400      f0�c ��̺��ο�J�}�[&��Z�@6oH+�hHb(�9D�?�x�F�� ~��G��#P�*ĔzR�q�23����6м�����p�Mn$��0^�a�R����&է��AF���-JE��X(�{����e���c�Z5��o���,L�|-F��R�&�:X��#P��3�+�)���Z���93)\c��PWK^R[��\6���gL�ח�
u�_�k�2�)�{�]XlxV61EB     400     110��eQf]v�������7N�;cn�g���c@u�	}~f5ѻ�4I�y[`�N{Ix��g�\��t���(��Ky�v-�=k\�I!�Ő�v�>����;y1`�F��������,,D8�~b���mJ�N胟8"�_5��et)R!~���c�\�/�k�V�d2�6��S2`���Ju�6���|�ˉݮB���}A�y�Nr>Hwb��GM~ytX�'�+|�<�@o�Ol�Dɉl*��m��٭�bp��x�i�!g���L\XlxV61EB     400     180� G�Z������QQ�`u�k]���m�����#����xQR��rbK:jFƇ���c@(��saN��2���F�`�s���/ 0lQ�:G9�DvF��j��j�,�#Ҽ֕Z�t!����%0X���/�Q<�E�k��\)!؆kZE���9���9&0s�E�Bx}�1���=IM[:�����TSW�����!��q��=ԉc��L���l\	���� �Ԯ�{U.�G��x#��"�Yg_�������j�֙���z"xD�E`���JX$Ͷ���4�j����2��Q�v=�b|�,�y,ݺ^9j��;��d���GЍ����RfBD��6�nI��a���A�p/<2J��$������*cs��XlxV61EB     400      e0�mX��L�~S�[2�K3�4��/��Zzhf϶�"��V߀Z3�!F��g�cW��`��0�g@��}�{�B�z�"e\`gbG���h݅�Z@�.���>\8�Z��:��b*쐳�.W$� z��M�o�s+ܔ�w�G�k�ԧ?�߱6�}���-/�Ҍ\j�ڇ^_q����ia��^��.�e�E�4�Ľ��fīE�R���xڗ�h�������!�Μ��:XlxV61EB     400     170��k�S5��l���s'qo��d׻D��<�	� �_skDڨb�e��z�֦���n֣2D����Rq^ђ4r��.	A=L�����ޖEL׎r�Dؘ�����iB�ٵ��>Q{������C(r�B�ɴ��%�QM��Y�?iF&�R"	�t�ۈ�V��`�ˆ���HhfG �.�[��gM���ܙ�g�V�Y�۴`-ޅ;PP�\�%��C~�kJ���&���݋�ݚ�ƕ6��>0R������4|O<�:�Ir�����9��L��p��J��c��/�'�*r��vˣr�4nT�$����lH�tMv����k���5�}qh������Ol���>3@h6���XlxV61EB     400     110=����Їq�����]��!�yY���԰��D������q	5��{-�*5�H��}%��=�xI:·a�����[���[-�~��;��W	/�GdV$���/�`ơh�Q�G���BZ��ɼ�
���$7�h�G��1*S8���ݺ�s?���Ƈ��S%��� �L%N��+�9z亖$���N�˒\�>]��Q�d��<~�K�6��F����p���6�s��յHyva�Ԧk�t�-*����u�V���w�u�XlxV61EB     400     140lttl�v��EF~�(��'�ˑX���FU����h�P�Xm[�.�{��!�����X˻�2N?�j#;�->\pi��p�B?&�aQ��ۍ9������΅��`$�����O� z�T�����RG?�`nv(q ��g{��CT��8��?b[��E\;o�%�W茪J�s����`�l����_Bf���h]ś�ٛ��p���ḡ�+~G�i�@D��|k��A'"�b
��/�66�i:�W�BW�W�]������i*��k�+�[���e�X}:����(>��5�B��چ}�I��ɏ�pg�>��c ��d�� ?�XlxV61EB     400     150�% ��Eڽ$J�O@�G�0ٛw�c��{�[ޡ|+c�eD��(4��Nb�x���+�U��>s��W�Q/{�(��W���/�=FAN���"����v���h
�ϖ����jN�w�i�ux�9�``���2���Ǟ��؊5J�h�66�3�U�!(I�>��X��9�dm����bjGw-��̊�}h��$�o8��n�w6���VIq����$]�V�Mf>>�H�D@#J��i�,�8�uݓ������&�>�]�Qыd-g�7J,�n��{G�x��M`���{Q?��Ro�W=��N�+#[�m��g.P���7ÕXlxV61EB     400     170W
|9T`]]�K_$�b�D���im�5I�RY��O�q/%�A�)R O���j��`���D��14��P�"O�!"�ԋ��E��	��(�xs��2�o깡���G��U¸��}z~=�x��з!��:�AW
��5�fbK��g�M�Zie��Lϒ;�ao$ŭ��8;ɓM�J'I�p���x��d8X%7ї�q��ii��QA��kt�ޟ��&J��A�M�
��S^� ��5{<;������=b���A'�� �Sd�o��A�����5�4DJ�R�� zń�x�0E��ߎmOE+=��sn����..���V?[F�6x.�.��-���`_�q��Q����~U�XlxV61EB     3a5     190��~r�VrG=ͧ��?��)@���I�\Ѫ7z�:�d]:q=}a)�ű�y��4�S��Ǫ��K���DS���w9/E��R�_�H|��L�8��UIRՎM�V��hSu5�þ�ej×@�j�8Y�HZ	�����B�M�1Δ���!�4j��C�Kz�t�L�5�E�(��&�{�jw�EL�T�/��~ڲ�WE��"ƽ����瘠?}\{Y�?Q_��X��י�\�5��Ɛ��nz�Z��ak��p�i8ƹӴ`��'yu�,w��b	,�nmڹs�b�"�9��=偌)��?��4�PZ��G4��˙]��a�(�[^8*@�y�a��)�kuru����;n����<=��c���Gk}�S;���u�J!�tޱ�1�"6l&/E.�b�C$h�J��