XlxV61EB     400     150=,�{��$�!��(Vj��q�|~�P_�:�l��YPU��3�Gpzh0PyC<i#V��HI����"SzMвz6�����Q��Y褅����+m�����]6�N�Xy��=ہ��b�]�Ya���N闘N���f%�,u�a���M
����&����	l5���R4��m����U�|+�u(�l��x�!H�9(�+9��8e�l�]N��o7�T��=�� �����"�h��آF|z#�)-�8 ��F�(�5F@-�˸��M�{l�_&m��k��6�:֭����s�7پ��O��*��}�
�M
P���3�@ �r-<D� XlxV61EB     400     180���9#����z��Ic�Nm��p$Z�<ݬ֊�h��q�k8�Ox������2l3rAI�z�v7�'8�0;�6M�zJ���Vu��.�1Ę}*j��}]$�Tg��(��Z�5�W���-c�:�S��Hf���cъr���"p�{y �+��A��W| ~
0��%�d&[� ˍab�)��6rn������a_�P'J-$�<'|o��>�'zV�y� ���v?�\��L\�ʾ�rq�ϸڭq.���d�k���U���O~�S��M
z��F�)�DZ�1�T��W3Fʭ�����ʍ�<�?�s���,tfo�zQ��Җˉ�տ�����c�p;1,�?�y�6
bq;2��ʥ"���;w��!ΤY���XlxV61EB     400     1a0�!M)í�A=x�����~�
D��+e5T��{��u����.�)+|d���RCf��{�>��'�^)�A��)k~'�1)���;땵�`�6���Ơt�U*{���-�h��nCQ>	z4��.&�����W��fK�;�P�oiK
���n�і��/_������S:S��wÕ��uj�'�N��x�yE�s5l�2)���4A�m)�r����{�l� A�G����oNN}C����AH�,���B7[��O���S��?,��"��Ӥ
�-es㑁<E���Q�����fx[A���<8�[T�%#qq�r�/��d~��E7D�;'��x��
��\���>Dl�)c K�3RȐ/s�q���H�����ebd)��17�ں����_0���H��Ϊu����HXlxV61EB     400     190	�uM<�Z�v���c-�j�9pBv*�|�������&�����&�iV(������ɻ�n�'J�k����'���uA>R(�~y�{,x]B�Ac���s�lS��:C�iK�n��g���K9ZG��0�V�3*�/�0g���Y|��
�e��1�	���ڗ�Z�p5H8&��xXd��¯�_o�; ��2�B�H�<:�Y/q)A5H�s����NƛP���O��O�/�J\�~GJ�G��Ō��;�1�t_��#(JVP�L�u����yn�����t\W&}��Bg�,��&�(���l�.[wXYjj!��0���Z-����	6'� Pi36ٿ["?���;��2h�ws�xW�}��)M�0�L��տ �ŻB7��a��#(�s�ߥ6�!��XlxV61EB     400     1a0����b7����s�*D��G�����h�O�ƞ �u�Zh�Y���8w�Sʹ��/�6��e���d����@���f����l�'�4�mAFZPb�Y1�)J/��jA��XM�Z|��.uv�U�{U��y\�����Χ�%j}�w6K�E��D��ț��g�;�a���5R�<]�]Crj��gv`�_��d$��(�a��*1���i ;i�n�u�_z�&�${߼'��I�Rf#¬��ɹqY�A	��/eK�	'��~y��U�
Y�x[>�_��T�l���l�׾��H>�u�-X[�o�;�r��}���ɭT`�M��H �h��⧀n�}#sc�6��~Id����r��:%�'4}��v�Y�{o��=���!�8s��}�#�c�|4�i�%��{#�J4�n���^XlxV61EB     400     1b0��J~p���5}/�n���5�"�Lz���!���&�)9�di�ˇZ��(�w�E�{k�z'�LӲ\�����h��ۿ��p�3����	�/�ߩ!�궟��m����t�B�>)3��썺b�ֳ�ㅙ�K%U=%��;�ߘ�å'�@���֗���;]uG$q<x�{���p0�ǅQ�V����U�"�|���B���x�p���-���ױO�q��OV��v��r���?X����	��q���1�Z���Y?pc#��u�P%E^sQ�
=V([@�b����)MR��KN8��9w�,�=n	��x�N�j�O��YĽ�;Nq�?��`���ږ�'�ػ��G�d	T���,j�A*���{�U�wS���TPB��>����f����X�����t�K>J��Cn�2�ď�n+~Vhxsy�Մ�4�XlxV61EB     400     150��l�(�ې9�q|��U3U�L��ɸ;u\NQ�"3Z+�w�U����4r�q�;�i�.��Tk ~]*���Х�0���1��;�: �V�vs�7�<C�d�{���;��?נ�"]�i,&K/4$�K�9��
(1q�l�B�h �CZ�-f��,t�%sD�A\m��"�?�s��֬�'�,��6��z��U�-�	�����5�ۚ|a���EK�z���Z�sX�3�{�X%���G�a�
�M�6O��;��t9����R�t{�@%9��2,N_�$��L�8�K��q�,ŊJi��ڝ�4��b� �h����Q���XlxV61EB     400     180�ء��i�1�"0�oY��!���f6/�����D�+��$�0�3��^؊\A����� 2��T���P�=�0�?�9�*��}Ď8��V<��$9��t������7О9�:AC�EB~����V�Fw�+4}<f_z�X$�Lio"��$�J��72Zt��?5IF�V󙴾�Q��JAa���6U߄���@=n��4�e�ų�#ʓByera '汫��:�~s���G���e��:��%P�p("J��$7��������n�b�Ώ��n�YU�V�6/�+5t��*�z#5�=m��6y/���V���S/
�7�k�P
EFT�Խ�-�\�gvF�fv��AZ�R1�Y2wM�L=K������x�^�Ҡ!zm�����V?D-XlxV61EB     400     140���iNߪ�.#�E��Z���h��RN`����z���a���L{�X�v���W	oV�3�+�u?
=��m!�^�n��R�y����ntg˹�ѓ}�J9�U5��5�9&P��Sy�e������������>�Oziә&=�
�|�9%����פ;�D�O	�WS�:J�,��%�K�,�t�ZU���!�l�� �b��PN(�i)���z��)4��h����ۿ�΃wm�.4m̫E����y���r����) �׏.H� \��$��� u##��m� %�����]��8k��5t<
���B�m�<�H<��W��XlxV61EB     400     1a0��Q�x �d�nN���w�>���h,���o�6��ع�m��Ew��V�$GЛ�Pe��^FT��9py��)�QH%�y�^d�S��z�j�2 �:  o��pB��Z��R�RG��㼴��x� ���p����]��zL����U��sq�O�E������QuA�f����w�O!�߆������1,=ߥ6�&$�ω?�6,:���<��k������fo������jd���&�3��L��:����0yo]���M_�x�� %[�<��? �ճ�5��@����\Td��
��["��e۴m�Ƭ�"FY*� S+J]	�A�.��筄�X��>X��P�ǔ��@�XaRbt�	`��gԡ��)�G�p��n��[h?�V����	��Z���G�>���XlxV61EB     400     190��%�����WCg���8�h�P@�)���)K`����A���%%�����ߢ�i*�4skl�I�Ǳ��H@���R
o������A�vs�׸�5|Hhݓ�6{i��1�>�E]>Y��s-�n�y��ΆI��;_sH؋�����3���\�ZlR� ��5<3"Z%�筀�HG=>�*pm� C�9
EcfA ��Dn�T/�x"�2`"�t(��#뒢C�&���Ce��vp_+HB� �x���z!�P;Ս�e9{L��d����TJ{b��0d%�J�2]�7����p�o�9�ףR�F�ʥ��ȓ���֢�����k�J��E�N�a���x]+�t�f��Z3�+��~ݨ�G"�FڤV.��� ;��2�������p�%���XlxV61EB     400     140�· V�?X���}�=~�Hy�ǜQ�P�X
s��\��.��q���n��:�e��Է�q4�>=}2x�90��˦��µ�&h�s�nv���$�Т/��C��*��Ic�X�v��T���3�o���B�#8Mi'���>��{��Q9w7z��#o�eI<����6����+CS<Ά�ڝ8�ir+ׁ�Yb&QG�8ٓ���q�.��1����-�>��;sBrCFtB�7��}p3��x�S��)��hz8ƕ|&n����[=�cҹ��!�E���{�ur�۴�x�B�zOc6���h�v5��43�8�\4bCPIa��6�XlxV61EB     400     1d0�;�n4"=�=FD95UE�O��@��� ���e�}�ݭ)D,�Y��c�U	q�N2�}h�A�����}�&c���R'XM�5�P?�@�+�Ý��ߩ�n�M�Yn���*���K�1�V�QK�D�>Q޷UW*���RE�+Q��}�S��s�(�����#�Tf	��kc8WX_��{(� �P#���a�ywa�l����F��G)�x!��0"2�n�`�a%���K�K���ڼpm�:;�+�N��? 'Q�݇������2�?Ɓ	NE�q�;�_髿-4TgV�]{��n��]�����Z�γd ���H�cl�O���;+HW߰2d_I�p�̦wF�P *l�?�����3n��S`XYQ����ЭZv� �;hb �1���X7�E�7kJ�-��#��gS� R��oӮ�P�}�ZB�.���5W���s��?�zXlxV61EB     400     170�+1�PÃ����@%ot����o��J�U5m�L��.��3�����Gx�e=���A?Β�fv 8�����|:��YO%i��=ŗ��Ro�ۻ�?k��4E�4nu�������x����p�|��'"����0@�S~B�KЭkج9��Gk�#%�fT��oc�	�%S��L���~�Xo:�C9��#D������SЬB�v�EZ.�����R焂�������c�W��\�^�������������`U��og��kʫɌ�z�p+Y����q�RX��ה�qV�܌���T,�Ȃ�I
�i�C������������3֍'4I�*�%�X������mG�ܞ�g��j�����XlxV61EB      c6      90"�P2��,����>o]H�����-�p���၊��;c2H�n���س��V�1@��;)�c)����޸!m*-حW��fcjLi=$0�])��BJ�&SV0�l��<r��
;�K֣f�tM;2��񼆢��/<�