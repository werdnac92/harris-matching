XlxV61EB     400     130��M��p�
���kG	ƛc�r��j�p�YO;���AĜ�/���%|J��YH/]R��i�y���7�R�PrЪ)'�̬N��*w+���8����nVo$N��:Z�h�S^<�hg,"�b����7{�;�3p���lo ԋ�"�/���?�aA����+�����~��K}v��00e��Hw,,ک����.x�P�����*�;"�Հ>���	h�G��� �5�0F���CaG�E����XG&�����m��bΝ����X:t8s��k��z���G�p��Ձ7��AW���XlxV61EB     400     160���3ʱ� �Q�cMsĠ\�j�#_I�FZف��vќ�i�Uk5�.�A�Q=#�@(�;{!��@e��?��D�N��w%��25�=6����3������8���
�SYM�������U\���}��^TK!^ą�C�-l��5w��t�!�/\g���V�%�X8����[/fRI���s����0O�����1I�F��F�Sܚ����2{����_���}m����mP���nuP@h�!#=�{��+�
�{_b//�[�̠�X����԰7��r���R�k��+0��\��M�{P���bӘѪ
���G�q)̸�"(3��vd��3-蘟t�ٶZ1XlxV61EB     400     120a���~���R����������ׯf�u0���\!�11��_|��i����G2qK��nhΣ�>7��)�����U�kp�Xvv��>�ߤa�"B�p@D'[��U�83��yN��%`��z�ߨ�K������R6��9/����>Ĩ��q�dBЧ%ʳ�K\��TG=E�Ŧ�!����՗o��c�9��p؍e�7���u��:됦�л�P,6��ϭd2>����Il��}��-z����p$m8ښ����^��c<@�R�.x�F�j %�;*XlxV61EB     400      e0=�K*�R3/��*T�(��|�.GR�mMgPi��%p�����xidn����K����)�k���v������?熰�R]��:�a�u Ϣ^�s�$�9���o�o��SW���=����xP������>[pR��c������F$xex\L��5�=t������S�q�_�+�w���m��2�o�-�k#�
�q����pB�NW!��Y�9��w���Clg���>�8?�T�fXlxV61EB     400     140`-N<#!���<��{�WE����P��5T�Ȣ���I������7������8��OhGl^zבᒮ���Bw�'kl�J��.��o��ka��[��J��j8b7��
:^�I(��0q���PBB�o%��%+F��`�f��㪁�!��QX�*��|
 .�:�#�ϐL�8L�k����Lo�Dm�l#S��S��3Z���{)]n��_5ih�H4��x@�H��M��Z�#����?��uL�_u}[T�Qg����|0`��M�V�N�n�h=��dձ�P)2sQǳ0��y�	D�iag��Yui�!%�ϫj��7,���6��#XlxV61EB     400     130��煯!��4��[.�O�~R��ٻQPM��!��2_�g�GT6`���G�9�;a�R�S�6�k�*��
���sA��Y���Zb
�[����ֵ2���> ��9���W�IT0tU�Ή�EhW�u�^� h���6�p����q@��oy���	)�;�~�-\���qns�����y?�h�?M�,8�︠��_~Z�4V���=�	�p�Ji�`E�@�:i�6BL+@l<l5���d�	��:����;�$R �ѡ/�m;������%\]���KFQHRz��=�2�緫�Ҙ���k��k��XlxV61EB     400     110��1�e�^�d�Ϭ��X�?�0x�:���1�x\�q�J��}�.�{;`��(���,"hPA'�/�M.E�
=�1�����9�؃���Pr����ɊG�T+�"�E�G�UGCJ"U^�W���YD�dc��y�	R������ �`�m�S�iMz�&vO���>�F�5"o��7���y��!Hth�a�yI��!��V�7(�8'Υ�Vs�(�m<�`٥��j���QhPx'��Bޥ�%�oWړ:^b���B�f�@�]H�KEJXlxV61EB     400     140������ܝ��L5�R����넕��b��54�/d���H�t���U5���a&�7S]��+M9�/rK=����e'�q��[��n���,q�����}ыX��n��]ط�$7�n�����=�������;�.��!=I�������C�?.� �z��-�q"vJ-�Q��sFf�h���=�^L�2�X��x-�Ћ�X�����Kg��b�XL�q\�I���R?ئ��Z��%�sg�y9���q�����������Z7����%����+vQ)	�r`��o�FЦ�W
�b|�(���ٛ�w����L���z�;��C3�&�y�+XlxV61EB     400     180Db��>���턗̗ey�8��f@��Ά% .�Gځ����j\��(X�;��2v�H`�:�(k��ۧe(2��{&�<�Z�I7+�4|��VM=BNoۡ�cm����Rft�ث��1#�Ͷ"c75�AX������#o#���O��(�PL�1ގ\���]�WЈ���j�N��C���[��H��l'R�}�*�� ��V��|������t����؉��u��C-l���E�\��I��6�� !�YODOw{�8:ђy_+��/��0������~�y��Q%ͧ$�2��M�p�ܖ#��	�
�qA�թ�)
���H�97�_�8���Y�Dˠ�r]� ����b�u8R��;��R�/w2�}ۀ��XlxV61EB     400     110����ZH��l�_�ʩ�SR)�Y	1ɞc�y����ٶ'�~DEE�?�nn
<�Z:��_���1d뇰z�ջ-�1�נ�h�ld���Booz��fc<"�tA�1�x���\(K2�.!�]�"5k{aN��P�SqR�=�_��6�,PH�<<�=8>�(A?�W]���dl�N���+��L��H�s6�ȯ�t$=~�����߰�5�i@zXt�%&�!�oN��R����	���A�*-��dp�%|��[�����Ο08�=XlxV61EB     400     110B)%7������ɷ���ݐ��%�T9�w<��䎦��\��L�^ENS��+��*��G�#��%�����::�(tu<7�����w���T���D�Z��	i1�0˂�3D*`H��~~�!��%�����C�]|翩�$�^�>m�-���l�ς��rq`�����<��8ς�0�no�m)�{u������D�X�vJ�9�7�<�t�;z�D1�ȏcݮ�pT�t8Ѽ1���I._@e�E����̞���Zˤ�*Ao{�X�r�k�XlxV61EB     1a3      e0q�&�þ�M�� 
&�kgC6(1= /��A[j����|N!�.�P]����B���r��
@�24����� �}G�O��C� ,itÈ������/~VO�)��{�WB�����V`էD�H��S����G�%�ʦ��E��]g�X�nc�M(�'4���B�6��qc邙f�woo= z�۔������jw�o6�gZMQEr-qaF#X�ASW�