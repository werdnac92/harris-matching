XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190�����s�ҷH'�㗸�=�z��,���5�/��Y�N&�;��%1,HN�<��M:x?�0DBf�-�lN�ʇRq?r*ڐ���=њ�|�0�B�"X�;?>�m���8U�~"(vc�!b�Z���P�FF�o��(�\;�P�����~ց^���l�k_��{�Vw{�rq�+ޫ�?7��w7��Q�)j�<����;�fY[�/����c*�W�)�������ᓾ������C������Jk�9�>���Zۼa �&����b;�+�?3�nT��M`~r������s�E_9���ʂi�Z��uxߝ7Ğ�m��-d2�A^=6�a����i{K�	��W��x���2�<)X{��֟�%b?Wa� AՓ�Ґ���חɊ%E�r�8>�S�o��{XlxV61EB     400     140Y�*�E"� -�6��B�T杷��ҩMq4*�������UpU���]��W���K��G��O:.hdF�.��	4�/�	�;��a�8$�b���F)Fg�3���a��^�L@N��+cr�gE�[�����P�H��V�ͨ�h9� ȘQD���J��1(����ǡ(m=�p��֪!;3�
���J6��5�3�ʆj%�2b�q��9q��bױ��Î���=Vl�<*|�X.���_�AM/�V@"�tg�����y��LŪ:�$��FĿ��sIL�79�9Ju{��қW��_�[�H��XlxV61EB     400     120��~-����������sk������6�����>�f�'�Ō�t�
x(@q79]�~b�_�j�ᙳU�"�L2\�xV�L�C^P��KO��|	� ܭ��C��8i;�Ì�����0���yq��R��0P.�ч�~$d�)��\�uL/ꀾ��,m�n�F�L�ek'�
0��	�C6�ʎ�'�<������Sa���I���:���o�����Ni�2�����M}P�`۟����e_�M��K)�M�&��6����?�C�#��u�t��L��n���KN�XlxV61EB     400     130:�n��D��=H�.�Z�W᭎#+K�_��_	GSｧ�G(İ���	sN��F��nq������˖����\iy�fHųb4���]�oY=/N{6��y�
��-�=��*�N$�G��~�������u���:{�x:�����ϒ���Uo�Ar%��^����iO�&(�l��oL��c�.�#[�
_g���*(k,'+��r8[�q-�J�������
suqY�v��U�ۀ��diZI�Uܤ�!̽V]���P@ 6%P��w䫍y���Ϡ9��T�ય�}A��.���dZXlxV61EB     400     120r�<r��M�&��Ȓ�3ֈ\�J�8i��Y�LI��D�m��F����p��m���5;��;��Z��D_�GG�a��5oV����&O�_���5P��*�M��:*zx��^����e�uA����L뼶cJ�{�JeL[�ϋRo:#g�G)��f�{�'�p�Ҟ��i��)g����f�?MZ�#��Z�� ��z	'��>�UB�bb��I���N�����T7�c!,_��a�Oǚd$��'��,m�| �Ab6�(�	+��؟T���O%�XlxV61EB     400      f0O���_@O��Y��/T���װ5�R�ɳ���������@Y���[�0�\-�t��s6<:�︊���p/��K��_:my�	xz�G�Rⲡj��t�C����疨2"���� 4���rC�q,��\`���TٿO�!����}��tvϡ�o��/}��@�2�4"p�u��h\�f_���k�[j�~��lP���]�J�g��`$�GgBv�mN�T:^L+��h"W��JXlxV61EB     400     120��mWN;�ݰ\,XG��?�!�A��7�NoNӓ�F
���ٍl��E��j��B�8N��z�n������ �wg��@���j�dw2����s�����y�\G����z��
�k��]��P��l�Y���'qwǊzO��w�| =�`���;`���G�E�<M�ĝ#kp�+��D��Ӛ/솩3�^̈5�� I��Up�t:�nX���_�=_9���<�������y�C}Y�̾�Ҙ�VŎ�/,���c0���5��w���@՛O�����'�XlxV61EB     400     110
�*Rz��cڈ-���C�{{���U�ܯ8��]+Ծ�zs���E�������È�G��x��[�A����+� ��N��Sz��4}S��A�n�ˡ>*|�W�+��y)4Td���0���X������5�h��T\H>�xzL�c+n*
�~�y1��j��k`-�� �M��;��Ĭ�p�O�eOf�(;��͋��:�+�i�BHj�x�g�X��&0���cG�ni��8�����z^��3�~~���b�G�����i=]zEtמ���^�XlxV61EB     400     110E]�O��z�CGWʪ��6���`[B�+�9����������f���Q�!�DX�z���J9��a7��0��mh1K��稜�8x��FwUB���	c� �$_�Y+��������4fvY�6��U����x}7T�A��o�to���ػ$Ѹr^G�5�-"?KD���Q.V�s���N��(��Ew�i���c#��U>�(�w�>b�vԞ(D���9������'/�%W_���;H]��(���=�V�<�ڣ^����JL���~�t���h�XlxV61EB     400     100v!
vVPթݳ��9�,��TC@�|��᝶��;�!��>.�y��ܧ�9�}�~n������f�������t
/�]!i���@��B�D$�gf��c�N{e�rV��j�����o7�c��7�W������a�9!i�MՀ��!H5�j�Leo�$.��#T����)$���7�rD ��<8<.�x4��� �#��-n�x���ͥ�]K�.��U��Q�8���e���gB-�-G�h��Ĭ XlxV61EB     400     140�h뭋 h �E/܍8��g�쫲�	��7�8�&�c�l�)M�SO��ub�#�i�B��)*�Z7���mF `�ynɑ�eP�����˖�P[�.�*y��ُ��5��}<)��`�j�݉֎z���^��OO~i�D ��������~L(7	�=�-p6M
.pLR-�����Irh>Ď��C�iZ&���QmK ��ŉ���<Jf{�3����ԭ��X�Ł�1����'�L�ń,1҄� l���{g8�����tj��O���"���a�=��n`�D���s��.���<�����p{Pjˢk`XlxV61EB     400     190h#Zd��K�5��Ȏ�Ո\dx�T�[���Ŀ���"���޴A*�^x��Ҹ��!B���VH�Y�
¨�Eh�g���z���RD-��`"5�,�"1q�u��z��_���9ϭ��~��7�2_7���)Є���t ��g5-v�u��k�#M�������a�yF0;�1��a8�-./hʆ�X����G;�< ����ѰGX��qj�0�8hXދ���'%A꟬�r��K	6�ixJ����1�Ș�}���:c�ާ�rf\xa҈Paot'���p��X�▞������	��F] ��q]lZ����nȥ��+#�*Yt�	�*O�Q*u(�Z��	���8�r��	�>e��{���*Ӫ�Ʊ�bg�.�i�3N���XlxV61EB     400     140b��������=�ǽߌW��8S����Z�)W���M�Q���{�����䡻�����B0��{6�ز_nD�ve�Ѷd�����,���D�(Ab��b����;)�}vݍ�f�4��<�\nPv�:��,i�*V!��~o�VTc.��?�X���δ�����N������N��$�\��U#��̀���K��0I�Kc+�B�W��ܥ�K�Ð��y�#�qD�I�Ӑ{��gWB,:��Q �)�]����RXZ	����N���˰QY��֜��.�C�{5��lFށOWf�̪e�]+�x�#�4��4q�j�XlxV61EB     400     120*�>(W���p��#\yg��{��`�lm����dR9W�)!�v�U�'�@q캵T��-��s4�8D6X2pS?�"E�Y��x�~b"�IS����T��Edsf"T"���2�o��I��]/-Z�E,�CU��a�|����r�O�e� ��@us�h�H&�C�o�8&oj��IY�礖ڃM���S�T�F~ݡ��<M����ԥ�Y{1����>5��z�۱ø�J{��K�6_�Z�����%�%C��$�"�u'�����uӫ'�|�w�)�	�]M�8;�~VXlxV61EB     400     110�W�໻��ۛ`����3�A���V���
�|����]�؜�k�	�֣�&����0���wY�ys�O�V}�.��]E��;��,gO���M:!�U�*����[��#)��. �L�=[nֲ��o�MW��Ϸ����4S iԥ o������p����L(pq�&>'xV�PʒM%�=�4;���P���hǸq���;oM��ŨD��,:s��,'r�he���PԻ�)Xͦ��L�D ���e��btSV�)7�$fTx�XlxV61EB     400      c0̊*e��G]`U�JK&C(��J�k8m��y �8����邻Tז��N��G�YGYTyQ�sӽ��Ѥ���%����5�E��k�"k=^�3t�
���~*���{/)��N`�%N; �{d+J�#�4�D}���Ƹ�H��7=,�9��m� =&`���4*1��=�R1���H�V�5]vh��v�XlxV61EB     400      f0Gk���o�DF9����UԀ��^�8�g&m�<�`}4�6�`*������}	��`�F!\�ܺw��2���)����@k8�'���5ξ�£�,�Ju�j�c"ﺋ�u�r�e���3�z���I�X�pS����*p����0~u���@x6M	�o�8��te���{���B��O��@�ijo�V�n�����]��!(�������[����c�ht�O��2���XlxV61EB     400      e0�VH�������M@/3/�D^{���}����|r�'��~�l8͐�&��[&c�_=���jW�>{���{{:Sw@h��\}N}dK��q��⍌+A��>��%Cڨ���-1~�y�uC�A�)��O`8X���=���}���I_3WA�&�۽ڭiN��ѳ��DyT~����FI��Y�8�u�C�Q��yg��m���'�N$c=���d�XlxV61EB     400     1b0�ȹ!�nHR�N�Ý��sc'��$\����ᤱ�s����4g�TB���-����`Is��\)��J�G�0>cZ�I�2�����mZSB1�#^�P�D��Pj0��r(V�L��;yiy�H����%��j�_H?nz��|�ހݢ��@���,�>`�B{�;&/�(�q�k���ŗ�;�E��GXN���ȭc4[m�,�.�@V<F�Ӵ_IZ�E�3�~�
?�GWVh�u�5�H8��� �u<x����(W�7��tG�>e���	L��d������4�#�^�L�AK]�8�_c"nhc�A<1&R�L2*��n�~o�qc)ipt.g��#�4�N6����o�-�h|�e x{�Ȗ��8Ga7�� ;[������{�O#��0����0���ok,����R��s��B ����P˫�.:U��XlxV61EB     400      f0��3�Jg�O��T�K�z�~>@/��SWDv|� �d��w��~�tQn6b�:f�ǩ� ��R`�r�*��<��*/��M�J����\�"(J������)�M���cLÝ#Q��QD�gz!�OwV�^ݼ�K�� ��9�A'"��O�w�����vTb�X�uu6N���J{��_Z- Փ49۪�q�_.t�Fz�ޒI_�F�������i����0$&v��qox�3�?~JkXlxV61EB     400     100L_םBu��C��Tꌥ�I�4��e��/�=��qȞ�)P0�>�۩�no3W�rv_��+�1ֶ<��m�J�IE[��X��j�.1���oEV�[���q�2om.5g�U�Ț��w2��C�ߑՍ�Q�c��m��dA��|cK�=[�kA�H��I3=ǡ5�"����_xN@�q1s6���D��zQ����z�3��t�>�����ݟ.�#|��Q1�h��mH�F��)^"����B��P��?���g��XlxV61EB     400     170���Tk��^ ����n���Iϼj���F� T��vs�c������J�X�e�_�J"K\�D������ ����1 �.�@X��L��0K�Ce��U�FV5f�&��b'�h�j#C�`�Q���tk����	B��Q㰸���0�>�����4�Ulp��.L���/e�f�Z�կq�c�:�LI~�}2E2!��e��L�Y���Z�R�:��L^��w[�mXt��_�4Q�b��z�i�Eh)T������;O���w�m�r/}w�d���<�'^{�gt�V���|'
ʙ��p��.
�So�����Q��9%����.���8�m�멌jO_Q�ɞ-����y����>}��XlxV61EB     400      f0��|�.վ,��C�5�i#)vK�V�'2e������8�q7au��L�l�Rr�\͵Nͽ�q3EA�YO���\����I)�^l w@��i�+0���u�YO�_�]�.�[r�Y��ݴW	Wl_�?�v�@��)-K��m��`���a��::���znN�DM�+]��h0I8g����)�I�"��yg��_���\Ù_v#y�B"��)FD�8 <�(��X�!f��>:�	ͥXlxV61EB     400     110ƭ�]D�/�E�����q& ߥ���Vo�5��]��	Dj��N�f���k(�1Z
v���1��+������	e�ڻ�������H�����:9��t�#H�r���Ϋц�~%��������^Q"����������T@������֡lF�� ��&m�yJy�e���UG���@A��7�Y4&naI��7���˒��
�m�I�c��-�#�F�@yq�y�2����z/��k�74����޳�f�[��0 ���o�@M�)�ÇP�XlxV61EB     400     1309F&P�诞>� �D�� Q�P����?���z�2���_�]Ҁ�!a��>}"X�qI�a�� �'��8����5,�qL���<;�� ��6�����#>�AJ*W9	��Z�S�@�l�J��G#`_z9c��Q��vV>J�s/�l��g��H�^�:��h�.#3���M*[��f!�=�%D�^ۙ��e���Dʌ�=�5�)��{��a�a���:y�F���%��	%��D���{��2,"����񲹑Y[��[hl'��K�Iˁ����-v/�J�l�V���������;ˬ]/XlxV61EB     400     150AS]G`�j�O��S2.le(`"�=���,�2����T(^��$t"�W�'zPG�p8�7�D��GGm�/��{P�[�Ԭ<�1�/�`�lUvm�U�*�~H��dṱ��x/��Ǿu�*��&�3�c؆4�!�̢���R�Z�LoC�f��Mp�}j�V�
�!�70BWt]�\;���:�7�賦��ᅂ��{#-7'�AtJ�h�>��:�8�1M�SK���-~3�1E�Qk
l�a�rX1��-�;P[�
d��bs�n��*���P��8����s�ܹ!X<?�"�Y�2��7�q�9����t=R�� ��`�l�J�����֒���ʛXlxV61EB     400     170�$C�̓c��	�e�,ns�C���Ŧ�ݮ�\"%e���M�td�6JO��ሖmd�p��}OTY ��p,��.�1]��?I�>��+9
Z`XSc��k
�Y"�˛���*���Һ = t0�P�Ī8�p��������	��<�@��]L���Cby�U���l���ά�����hS�G73��z6��� ��ۧ�sl�1؇Cf̣vܐN�x�'���{���o������^��<Ze������V�:GJ�ȎC6�J�
�)U�&@�&9M�$O�!�%��_�ϖO�&��Jn�'}�}��8�3\��4l�0����q�۵70 _p�$}��X��Y�+�/�Q�G�����q�	�s�XlxV61EB     400     160b���dNxV`��;�uÛ�GE~��^�� ,�@�d��,@��a˶�p��F��m����6�׿>���Ѥ��>\��6�Vb%��2M��v�N�geU/G5�nu�%���8��W�tQ*�;W�/q��;7O|�T�� �5~~��O�3�K�%����`�<kI�s-�ʢ����l}�v�{jb�}����H���� '�M�2�C>�H��w��U8/l���
^n��U4J`��_o���"tx�C·S١�jK	�!k�%ᡯl^M�f�s]�qz�O��P ��"��ў�}V3��V�@��&��d	��(��L�0"YC7"U�(��E�(�Jkz���!,\��P�XlxV61EB     400     120)�bU��Ɗn�wvx����j�#3Eݡj5+r#C�#oi��L qt�s��^}8	�ǟ�7g�檓�_�*��,�l������q*�x-��ƟFq�Jmp��(,�ů��p%J;�E���M��:h{'ߖ|z�(�ٶ~+E�(^Tb�l;��Z�R/�[8��6S�a2Cѣ�[3XghN�������3:j�X���'�����4)Q9�x���@0db��jk0輣J�tc�?���&[H\0rｰ ػ�d��x��4���/P.�[ܼc�c`O,d\۵�iI�XlxV61EB     400      f0��"W��6�;9��،��O��M�X�q���N�r���)�����n*|�S����r��?mp�/���5^Ί�Z�\�5��sr54�{1'�%�7�E��)G��8��_2@=j��R�r���C�^I����1��������o�y�/,������e޹Ҋ*�E#�F�mK�
���Oj@�>�u�d�\I�?~ �U�d��KQ�N�����/?R��"nѣ-�]cS�/��XlxV61EB     400     150UG
��B�:j2��"!�\M��@|�e�����!��.Q��3�M��;T����'qu���E�	u|�!1)�~�Ŗݧ�k�K�l�F��>���0�BӨc��؆���.�c�w��Ҳ���'��x�	���`̑���¼G}�h��uK���S�t�a�MS�S���xW)=�6�ϝ���TjĺT8�sS��B���8�'h&u�$���J�=e�;l�H�ck�1	�����!�0���ӎ��R.=�����]���j��j�}\ˊ�����J8��Zь�/H���d$_�>WL�q]h��
���)F:��Z�B�� ?!��%g�S6�XlxV61EB     400     120���&�n��X�7�{��@h#���Ӫ�B���I��~Z��B��?Y�85v�~\�����>�S#�`?3�,F���h=�j/$�M�*tVgt�#�C����ߩ�b��O�,��!����\-��V �v\}���K ��<j���͹7�n�B���p�-���g��{�W�5k��R�a���6�$�{f6��� \C��Ӟ��kk�H@!�	c���j���D�1��o�Qn��e$��.Z��ʊ�� eUm?W|����$��=8-䉅����G~�!��-�pXlxV61EB     400     170k�Wr�R�4�m�%�#p���UTFgaE7����U=��5���n���Ha#��ǯ���ؒ&*��o/&�|*����zq���DP���zbՁF񹚁@D��sbH����z�*U :OУhf�4���gx���We����TQ��;�����iP�GU�atJ���#�`ͯ���9�S�`�=�W��u���#Q�b�?��R�Өs+m�����a�k�r��wV�>��4�u5��ܲ������o ��p���<��4�G ��bz@��5#1h���2*ђ��}�et9�=�BCn�PVXMD�ɴ����^>��3���s0!;;��,����f��h"9�3SX�e9 ]��O��=��E�XlxV61EB     400     160w�&�Ê�5��E��D5�y�0hb���d���;	K@;:C��� �п*�A%:��[��?��2�@���D+;�+��l㏷bC�7��7�;S+,P;���h �,.a�7%*�e(L\v��
��|��8t���D��3"�O�k�`g�|^<J�Tp{Dh�e1'$��ȸ#!w�QuC��N�J��0���G(YGIAO�� �������v9�V�����c4Oq�j��<��~�Z[z)	�]N��]�������Ű��x��AA�n:%qD��e=��&�Qge;�y���������`oHɾ��}]���(,6ji,�gX�1s�G04,#*�؃���TG���۳��XlxV61EB     400     180���~��j�La3rP���4�l���u�ߙNL����I��Z�j>h]�����9^����5��ߓ�8�,F�O"'[�5��j�70[��T��[+�1r)�dlix��4'c��o��S�Q#z�y�k��59��(
ry �N{�g�+�V]4ݜK��@{"�����i�ݸ@!#e��ť�'�f��*$u�4V�
������49
F���vvdY�=��z�H�WJ�4�K���4�D�!�c�/��P&���wE��t����=��R��e�����)���Q�3>�f��vޚ�Ɗx�iLcOQ'�[�����Gd�'}e�c%�ci���	5yv��9�A�QP|�iO�]-��[ ]��΃k�^�:����h��P�XlxV61EB     400     150�%Ҽ�Vs'�����!_��h�"h�Gq%�Ⱥ`��BU�^��o�$X���z3|ĥ��F*l�-�"���p��[�Ga/��(�'��1��#������p^��FK��ɸ!�n'μ�|�:M��wVܨI�ٙ csz�&0l#;L�q��c��\w�ez���Ȇ-2V#W�!?!�5����O S�[i�׭���Ab|����f�6�<���X���W��z`�� �� T��8N�;aNL�#�ͦa(��|J\m��&�]Qh�OX�ʔ	�H����D����~�}� ��qI�n����:�&}���z�Y��=Ċ��-I����P �XlxV61EB     400      e0�-N^p��xI�\Q�Ǜv)��/��QL��e���_��EdV�Aqr?2	K��ǂ��=�O�i�ry�@����$m��Ӽ�Ԥ� [�*��NsE$�ػ�ٴn�
��$�]��łd&��d�I�=�mq��(�����Le���]n�_G5)
�����*��)�(5[��=��1�!پC�������^s�2�\P��q,ڕ?�M�7Zc���o��e�N-8XlxV61EB     400      c0e[�5�����7����]mZ�eC���(����]��v6�M��M����P�@|��a��;������ +P5�����3]AE��+U/�׉�����4�G0�I9# ��<����yY�����r�t֙]Y�����z�s_��n/K�5�i&���p�����(ޥ��:I�#��`�%��K�W.�XlxV61EB     400      f0�@22��}���k	�$u�K)����?���^;)��:n�"�����3����l��ҶX�B��5���hI<�����!�cPj� �\P!����"���hQB�%�p.3�jf�/��j�^��=lrS�����.Q�t�\���t�+QƂ'��t���+��`T���fkw��Q~��A���²A�a�����М��Ym�LUX��s0�b!|=G�A�ٯ�M�HXlxV61EB     400     100�n�uET�nyf�N��D�`�9�T3��pH���H|p��h�t�B�Q��&Q�N�K�X��DG=� NtqD���]�����@Iv�aF��j���H�ǁ�~�F����2��5�G���S�?�7��6Հ�_A��QK2�\�r�(y��Q�8zV�����vzfl�%���6w�I��s��� 1��ƍ�.YR0�֐ǾW��0�`���)��s�w�<5����8� ��Fd��"�h0XS�2�=t��Q�B�g�6�;�)s�XlxV61EB     400      c0�w;4�����ps�s��P|G�i�S-"@	���F�AIŭ�4i�7����ͩ��۝ǋ�R��VaFW�a�y����\-C���
;���vf���3D  �"5�n�CHw�8�W�Wl"uT�Y	�f)�we�4�A��K� �:H�ƅ�}	\V�Ѡ,t��e[z?8��W���X@T6�U��#<"XlxV61EB     400     110~�{e[{'�r4��WyT6��i9WH�q�����Y�q0f5�K��$Nk��@HV=Þx)�J4E��z^�Љ�_����f�M�!�H� Hn��>�m����\��˻�f�K�s�Q�r'"X��0Ɩw%�hf|����щ�sq"&���,DѰ���r��t��ϡ}�0p���*�X�|}��r��o�G�q�/��"��rm��m3u:�aHc�c��?A���&�8���Z�[%칦5s�����-;�@�e�zN6�G�;���BXxXlxV61EB     400     100�"}�σGK��ʟQ'{&��wY�M�Q�ﲐy'��w3q8�[�����G҆jr��l;�~f��v��m��qH��샠����>�V��w�U��3*�rS6] ��������J�=���=_����$�����,��wlTSsM����UQS�?b�!��
	�9p�{դ�Aگ���ԍ���%��姃���W8__��9�TQ+�"�q���:�{M
�����p���m^��0�v�����E3�J\XlxV61EB     400     140��������G�MRW��Ϟ����o�0��>۴�k6��'�Tݸwz줿��c�m��"m)F� >v��u`l��0��\�1i?�3V����*=T�Bc��	���-�`��>;ZS?�0���K�p��z�Fj�6��1����dX����s�ase)6p�C���/������_r˄��	{�����#F����v�U�P]�c�
0I��_e2��n㵟���n�/=cO1Ҕk.n�-�.��m��C�F/п��7��y�)S�Me:�B��M1�8ȍ�@�踏wޯΞ-���z�(�>���|�����XlxV61EB     400     1a0��`��� ��F�3Z���Ocq-�o˾��f�<�U�
�6o�3��|��_�v�Ԓ����~L4;���*�R���L`�|���4x5��0�P�|�+�0��"�����������9r�z;Z�����(�^̏��!vYe����e���K�����ã�m;��ͭ��鑴_�md�Ҳ��_%�DW�G���(�Ogw1 �9��V�y�ux��J�(��soΟ!Rm�m���[W:��w�A�5l��_��	ۊU��X�`��@�[��w�m;�F&����;�R��|2skuN�kYUZ�F[IG�YQR6��"{�h����F��7�~.�q ������J%�r���r�ˀMӸ�|����Bi��'4�1S`KZf�n�Lqw���J�_
@����-��X��v�U�XlxV61EB     400     180%*�~d����X��q�H��ݝ��\p���ö�d���Bcg�u�,`V�C W+���X�����G��P��}�� �;�'��)\-�2�U�l$j�1���gvU��z�K>f�����ӹvX�ၕ[v^5�b�_!q
^��1ľy};�����?�-�N,���߉9����E��g�:h�O�>�7ঈ"ǯN�S�'kM�S�V����ؾ#��]��e�J4�T�ۡ'�=
4VO~2�kD�S�w>���f�D�d<�(���r�=�rx���:Z1C�\y�5��gh���K���=�ȔTK��c��sr�Feɓ"1_�-��t�"-�;���W��5"��V
&MЮk21M5��1���C����3��4�cuY�	mpF��XlxV61EB     400     110� ��	,��⊧,4U ��q*ک0S �ٟ$�}�Մ}ea��\(ص�@��q	uI6�˯��+�ĺh#����y� \��;d^L�d��'��ru�Ԁ���f�����Wx��YrE�jz��4�O�X� 8��}X�C$��1�����9�?������:$xA��\�%('��%_�7p��TWj�E�ND��ृ��4����X�h�ʊ�WDF�g��?#q��O��z!ށy�Ϸ�=n�f-5 ��Ww-�r���Y��kƋ�cXlxV61EB     400     180*�\��TX�Ӷ�Kx��4&����Eь�?��rt��������񁄐�a�g����Xa���1��ߺҳ!�.�����F�9�
�X�Wn��$�˄9����
T�ܠT`�Z�F����8]�?j:C��D��,z��!��-� /�'),��B�^�  ��AL���h󽄡�Q��-�v^��/��â����2Z2�,7��<��v[�-�o/���,�64��ϻ����H`���m��~!���D��F4�8t�������}��χ]π�,�+�:��X{E,މ��82Vq�C�!ñ~�[�$����C;R�1w��w�0(�^�Z���x��{��(_;4�ϣ��wh!�j���:�u|̣����XNWXlxV61EB     400     170�[�Z������B�TS�����g��܌*�������ë++�Z���<�����Z	�`eXvhtL��bOrM���7�G�T��VğH��ȡ谚�K���godi9�M�pAK�[�^�����E%�_�2!7\�Ѭ�&��8Y���/^/P�׼4�H�o�] A�J.Y�إ�y��i)�*��'Iw.� �����R��|�j*�0ƮÓ�q�)��6EI�,x,7�>�c(� L��.��6�u*OBXF͏tdn�,��B��ʵS/� ƺbK�e���&�U?��T݃�!��x�!9�nQG!ۑ ]7&��ɤӏN��g��;��8E�@>�&Ar��XlxV61EB     400     140�`�;T�İCm���>݂���AXeM��'������-�1����0dQ��Yg���S-���879Dd���\�{g���}��뙐��+{�$�4��m��0D�g�"hM'!4b�e�i"����F���BS��[*ĕ���S����b��B�I�����ȯS���
��!K���	eC/���)h�����������(`iU��^T�C�p�e��l"yʴ]|8��rsҐ�����Ug2������m=!��=��;�-T�Mmc����)��tQWg�3��6#��<�8��]7�VQV�5{p}�/3�Q��XlxV61EB     400     140��㥛�_�B(n,�Y��t�E6g
�67����cvY����VS�e|Ƶ�}L�z�D@�,���[�W��uTw�q[�r/���n���K�v�0��Y�,�T%2#h���#�Ь�U��
��M`}����{+s�Z�p�]�k�8P��Ǜ���3PN��l�&�!����}h��X�r2�R�H�ɖ1�s[u듓Ňw�����C{�������U��F__
�DH���?�X�2ڗ�R����މSX��3��z4j����4��#1�
��ܪ¥�˛��$���%͔�2�O��fh>:�K�7XlxV61EB     400     130j���al>����o>�G���`��+� nZX_a��s�)�RG�N�Zh;�9qz�W�OTkp�}vK9���	h���p��%8H֕-�3��dƾ�U�Y��`�v1��ڙ*m	�3F!V���I�Pj�,�ɵ̬a)�\!����l�Ij��ߥ\���$/z�^MI�Mִ��F�z+���o�H#�ŧ��R����)��rE�W�*^���C�DB��������z�"1��4�<��.5�9n�b��ϮQؑ�����j���� ��h`�f������d,��K��K�&y�9��S���<a�?h8�%�XlxV61EB     400     170%����qR�p��d�`��i@�_{c�-b)%2��iD�9^�mw-wi� �`�;'���&% [��t׶4긤��}�/z�SĴ ���*??	�H��_���ܸ.U�>WH�U��|�m�\ᩮWtK��[��^�z�A�_9]Y��[Lz��א��֩(�@d��(�m�{C`e��`�c��W/e��lQ�S &.��z&�EϠ�O9[� Sq�찧/l�	RL.≨Q$G��N��b�3��^�K�N�m�6�i�y�ء��)�h��!�_�II�~]�?Mdb��#�p��[���R*�F>������Յ����XHC��ؘ�"��W��#o绌Ӭ���(]9��諾�I V�XlxV61EB     400     150HQZc��,���N��."�E�ɶ�;g7��c�N�?8��OV�^*8ҡ��t A#�DG'�BF�y�S7w^�M-�:�t·R�vb�P.ԯ�g~`c��{�u����ZW�����3�*�8k��q�ZtJ�Cg��S�{��A�A�B!I�.�8�o�u(��1G�>	�My;&`m� �q!� �O�����d����(Q�i�)�z��k/�)���C�}�Tz�\P[l=Z�Y_��+�\�6�o�2~��%K؄��~W3/:n����73���Q���/'�ռ�Y���vb��Z�l� �:Ƒe����B�b/Z��q�XlxV61EB     400     180�!8a�<����H	f��i*�[�N�h�m$��7L��x�O��S\p"���(�
\�O�tM_��=x�d�^�ِ�������jJ�C�!�*v*�#��w�jn����03I.v���Z�l�rS�M��(�x��A{���[g�-�T��j�i�Q�qT�zଦ<y��Q���n�9���D���&�O�) ����=���\JAO���R��=W��뢑N��Y�H̢ر�y�m�P�X="A��k6�ͦ�;�E37=��������u�W��|l��mc ��s� �wy�����G��/�X��b�Nz�h��'�Q�����@H�K"g�������y�C��[g�M�{�r�ZHbI���*�AP�q���U�XlxV61EB     400     180��� �x�\.K�P�=޺މK�ڛ��=�.���N���&3����6d_�� =�6Oa#��Z
$���l��#ɫ"�w�#�f�牢��I�1�Gr�~"k��^�`k�ĥ7Hw���@�����Z���~�B��荗�z�z!�IyW\ʙ�d�a�6�&e#�>�SG5�Ԗ�m�x�إ	��AY/��<g���DB͐����"5�"��؋\菖�^�lA�
���CxޏKO��S�� |r��X����A&CK$y�*v����/�Ň��2�ƻ�}�����v����3L x�Q�Љ�!������`6��ÃQy�@VL�H��G����x�d9I�x�\B왔y�K�Q>��h�8���s�LV�����XlxV61EB     400     190�i4�U����tc��d��y�.��X��e*�i�H�= ~�i�����9�� y��	q~e��K_	�b-~RmL6��vU�G��!�z]�=�Ŷ�������_�&�*�Ѣ�8p݋���λ8�`Z�o���5h�\��1����:%g���{k�b��W���[Ha(22�A]�w���u��[�n�^p�&G�:�i����L�N�*�S���:��p�ՇVec�Ŷq����~�pz���4k�������N5�2R�NzL�s6�]5"7�OP��N���ݷw�L�Qo�
�>i])Q%d�c�c6��h+�j�?ңXrK�{eD�M���FS���y��-�������*��۹�-�u͙.���n��3njRS��3��f��XlxV61EB     400     1b0M�.%��f���帀-M[ha,J_���J���in���4����Zc7Xךd)�� ��>�7O���~㾸w5�au�r�y���A�ty��ϱˇ64-s�p�j������L*�
h� g`rVƕ=���@�Kt�o�i�G�ʡG M$?6�!� s�'�A���y��	���0{���@*yz�alo:�z��Q�M�%%��~R�v���X��R?��#�b?^mrE#�n��#ꌼT�,~κױ�'GL�O��� ��������D�'i�P{^5�e�2�8���.�� ��|�?���&W�L�����OGp��;\9`l a��X�9^|�������M��u$�˸:�>Z��|9�#��	�@A\"�5d�{��u��`.��F:�ZTY�LLAz �-N*�4����дW8}F<���ʉ6�XlxV61EB     400     170����^3�n�yu ��k�?�3����1��хwH.���d ���;|���|v�NTV��tM�d7PtF����^����4�a����7�uzC"�|xr;2�>�LT����#��3�_;��"MXŹ��*X��w!�RaE�1m��GL+DL�s�72?Qgoe5q�KO}�`�bԴv���%� I=���:0���8O��3K۩�<�Zjy��Q�Zn��Q]8�%�gc0}w�i��E
�:����I��z���q��H�U|��8�|�\S4���6/Rp}�J?�I��~��<X�uq�
���a$t�ւ���X�Q́l���o?�eVn��ZX�ġ�G�kM8ެ���`��XlxV61EB     400     1c0��y�17��h�*���Hn���D�R�@�l'9ʷ�i�7����=�����X��I��C=�t0�-���&e�o@N�_��Or�~�$z���^�=!f�w�S>��N�� 4z���
�P	$Y��0�\	;C�K=`��A�9p߬�'����╘�k�� �iZ��i8�1T$'������	�a�A39�珩��xN���Ns3f���\�{
A�e�(�N�t�])�h�N��*���S��-���wUF�����5���t�l�"L����I���q���!��gW��A5�������+nɾ�Id|�Jd� O��;-��."�&!]
���K��Lj�K�����F�S�yC"�ߌ�H<�S�� w��8#�8Q���dFP��.���
`[׭e�YU�VI0�&��v>��\�>O���ؿ	J�D�0�	6��YXlxV61EB     400     120v��症��V��y���x�)M�L?x͗?���&�m�j7�(�Zl~x�Qc�`s��n!�}�U���6�Mf�='�_��327�[���z�;v�B���M�̧��C����b���*�F|{�;���4�WF�P��`5%A���V;�v���ږ>��Ӫ�fE���Z����� ��7¾3Y�E�������R�9��OXِ��T;�� tJ�x�^�?�u�;>_ts+�B�9���,�0�ۘb�l��=5X̻_^(�!�����ym� ���XlxV61EB     400     1d0w���R��ҳ�R���P���܀s���ͥh�����0�T��,�6c��ۘޝ(���$�- ?И8\�'���3~�ԫ�r=��t��$�k\�aC
���U���c�^,��J�֭��
�B:�x�H��nA)�*�o(�K���ݙ9;�ŤnUv[�еs�\,7��j�FK�]��<��n�d�$%��)�}�=W�S-�(��+%�RٟMuY�d����T;��_�&+��Ù鲻i܀Z��s#m���HbnM�	<~mn���Q~�|T
�$6�x3b��{�kTc�	{;�)e�k:zh�����*o�7>u����b�:�ϯY��\��NO�����"�����B
؜��RüGG"���xD`R{����a:ШYS٣6��������aY�\�h��,�u�Y�o=c��C�H���ݟ�H�������ί�<���M�E�Ui׮IF�XlxV61EB     400     190�*4*�m)��U7و?�����V���-E}�k�RG�&g� [	{���0��d�ަk{)���5+��*�ˏG�12�}�#��f����a��O�`+���t��[D��^"*���ń�,�zF;)�C�6<�H���b�gۍiΖ�?�	��Ɍ�N�~G[o����0��v#���勢u̬�iقԎ�L����=��.1ҋs�%ર
l2��8�AG6���`�ʧ�#�kKL^�e�G\0��9�d�G��E�N{�Rhd};`�,�g$�Z`Pԛ�w<B��X`D��!��CؽK��׽�KG���_>�����?哇���h�A)m�~���}�:	��5�uz�@_ɧku���|t�+���"m��=g�,��p�M�jXlxV61EB     400     1e0*o3:��
�KN�l��D;>:��F�Y�-S�Z��C!	;4�����G,���X9�l8��rR�z���0�2�T2V�7���������D#��_�o�gL�����f{�ؔo0'~<G��[�Y�������CN��p��U�V���.98�����8r�:@%��>u:���Eq9U�#p����tܗ<��'$~"l�����^��P��H�ބ弶��ɚd�_�J��.�}�(g� �1�61^zP�N��a���s�����`�q=|�r��c���*���M*�f��2��8�-]����zn,��pDl�$�j*]^�ݰ!�,i��>H5�W2ew���|�PjnI���fS����>�P2����FVA��
x�1nA������>��w�!G�^�-?W3����������4а�ƀP@�/��A�W�a�7aܙ�o,t� �D!�ƍ�O`P �V��3�O:�%$���x��l$i�XlxV61EB     400     150b5��U��_��r���Gc� �eP�UF�rI�ܱ����	��f)�U��a��j,ȩ�\�g8�r�c�ն�BbI�AT|����n���
�q�!�6�<����	D2�Orx�	X)�����[y���I��Bl��ˠ_7�C\�Quf�q�mo&>�֕o��k� �m{W�h��R��d�V�V�}OHx���� c�..��ͯ�,`��TR�2�*� Bov�f����P�l���|Sw���;f]7�U%сw�|����ң���)�
d�_b[��U��S��*��A�ּ�5�=
��N���iE����۰��a���6�߰�xXlxV61EB     400     1403��2v�A��x��~#d?��d���Ɨ�����\��V�&d&�;���t�q��ǵ�ۏ~���Wf}�B���S���� �ı�-�|F��ߦ�6��Z\�~��4��bW�Y�Ou!2����][ɸ+��iN��B��W���,�ߪn�T���VlN����#=��~�h6��^(���;�����<�l���^>�K���Hgk�5$�9o��/�~�浧6\6��'!"�w�㧁�D-�O��L�A��V�+R�R��᥹,�� QA�C/R���@>2<��Tl"ޖR��1P_m)��'Ȣ�w�)Q`c�XlxV61EB     400     1a0#DbB/䦞��82��:�!�T�m���h�����f�X�v�{Q���n���;o�ItSe��M%B{*<O������d��^�ə��'�s���-�ܣ/	�<6�M93�<���xx\�)O�9�vȈ_�������膂HI��|���S��,`��T���O-���Y�Dx�b=���r�M��M��p�md5d����}d�Y���␾a�v׳�T�ꇁH��OT|,ip+Ũ[:eAeX� �(��^���Q�y��j{&��t�Cx^�N��\+[�1����}�+����;����ɑ�p���o�aC�a�� ��-z�>�����\����ǀ(z�~���O{�B���@�W��j��Kfi�d�B�.�[Nh̛�G$נO�2���K?�~��"�l�3�jXlxV61EB     400     130Yt��T� kE:-�m;E;Z��'j_5��0�t1'"l��5_#G%�u�f;��]��h���ws�q�c,�6"��[H��E~�6�鱟��)�@�E�7��������pj��JW���Q�<���9��ȠW��ݑ�*K%�#���/#B86'��G�6��7���}�b  rS5��ZJ�]��qX7Q��*��S���(`k�J����a�5�BN��Q��bVL`]����HNo�&��X��)'��2���	���0�Sh6(����\W�.=���]�`]�dj;��yfR"���Z�XlxV61EB     400     130���|��b�����θ��sh���lX���ܥQ�����ͼT�m�r��!DY�S����'^I��I修������K-�BG��K�K�S�U֨������`����A���d�k��#4�2�7#>�̝�OxC!�3��B�N�����#�������wm̎x��ۍ8��5����2��\��2�~�k�n�R��Wݑ3�x�:� ��G�c��0[�W��y#�;��$�P��Ol�!0��E�X��zh� q���pⅿF%\��n�)=�ȌKbQ���XlxV61EB     400     140�q`.��#�V �+���T��
��AI��TG��⶘Π���A�ym�*Alf�q�� Q�t��͸������i�k��%o4�Gc�EV^
�F�Z�n�IF�Boj8X��瓶��̤³���j� *�*a�^`q�Öt��O��t;eU얫B�+����s���M%�މ8B�Y�RX��" �AE�AW[�Y����i�S�ķ)S4�1�/��c!V�^g^B�j�ٗ �w�Hmk~�-Nu!��r�(`��bP��5o=%���|!"��
�*����6S�>��y;_��|�� q��/� �	��| XlxV61EB     400     170�	c�n�v�ȃ�A�X*�sK�E�/MSw>^9	/sݕUB;9Ꞔ1�ʜ~b��{�HN1 �}�T���+OEE���ʯ�$uN��w��j��XS*7�\���"��]k��%��6
�$��9�]��M.��x#�[�)q�x)���鯬�e�@�G�5�W9O��$�O�*�vԉT��!n9���ţZn�;{�.;���; �����<.MO�u�_�(6����xY�|�[:;���8�Ap-�-�ʚ�*����-$���1��R��7;a�h^���]5R(�t�&í��p5��Íj�͙�	kW��������k���A�R=C�s� �-=��W�4���|�x�q�yVb{XlxV61EB     400     1c0��櫊�B$1�>eA�a	b���9h@�>n�����'��<��Z�M�����7��)��*�o�l0��O"X����K6&u@"Ћ8����>7�z�9�ݠ^�ı��R3�S�ā��}a�J�<�G��k>�x�68���wK�<	�����O��~;29X�H��*������t�I����H���މFW�e�=~����m�\|3�4�6�Thڶ4��K\���F�Ҝ 
ˢ�XBG�d�1��~����뀺��a]��2DB�7t{L�*�"�qpc/_�ɖi�u"����;h�L�%Av�cm�G�n������H-YC���/kГ��!N���QD��۝�̾eL���o���Kڴ�0����Q\�{Xns�\ �%�R{�D�*�w�'�ӺQ�����^����ɟ�m��)��Ĥ�l���*����ް�XlxV61EB     400     150Tq*��e$Im�w@�W8:�^r���G�	�O9+����}H���� "�BُM��Q���z�ꓱĐ")H�L^�&[�*(�n�N�jmT�߾����`���u�".����v*���,�~���%���;d�q
g����7�KB>O&�+i������l'�j!d�zצ{��H����,�G8t4�u%�Ԧ�<@5����6ȥ+n0���+����۰�n�ܙ�9��̭���$P)T��).3y��=6�e@�0ea�"���q&#6ږ�ɼJ�e��J�
�P�����;�f2�0�#���`X5ՏQ���G�8�G�U	l�,\β%pZXlxV61EB     400     1101!����<#C��eb�!WQ��2S��	ЭY��?d4�3o�^ơ;�,��|bK�0E�7�)<�;�(�7��E��׸���`�Ѯ�`��ZQ��Z�PU��DC�xy�=�XW4�
���?��ki>�M���<
�IS\�����nPQ���k۞�V��(�8xs2����Q���T�����t�v���Y����,���!�w]>@�jJ���:G1��0�<�ɓ��M��ò4��48W<��S%�w��.Iy�r��t�(��)q�
XlxV61EB     221      f09E����҉�&��@e5��czDuՏ�CZMI-�Vq2S����Dw�^K���zaC,��;���	,�;J���@H�ѽ0t�D�A� {�(R�8�l�7�ē�p�f�z�o̰�mSd�_�lz,��NB��Kݲj�{��9�TM�#��`��V��}2�P��!���Y�߱_Ӻm$�4��!q��{��0�P��	،}U]A8�Ϥ"���g���-��)#���;[L}����\��l��