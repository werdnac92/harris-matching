XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     1a0_�?ܓ�|Yۘ�>�L*qj��t�0�PO���yvr�Ԡ�|�e鐊�vd��4�W�/�Z��T?��^�!Gr�{��ȊE��|���C\�q��u��٠���=8�f|"���M�I6/I�P$��1Ի^�Żugp
��:��g?��d��qԇ�CI�c?��Ũ+����S�@=�lw�3�Y4(2�˟h�y��x��(�;��A��癱�d�-#�*�ܝ�pq��d
�����t�I�4d|Z�V�<�Z[���5�v;����U
�ICx�;X3#]z�����������g����A��c�W�k�޸�����|g�8�����U��67���Q��BHǓC�f6t��1��)��$*L��2�>;�?�!xW��K�k�S���$������3-�zx�ïK��컥�s�XlxV61EB     400     1a0P��_����ї��~l�Pa3���+��l�*�<S��&N@���s}k�Y�`��z�/=v%���
�[JN,�S+��>��!{�ک(O|}�˚��~Qω�礁I�����La���:��W9e�g����8%L4Q��Yt{g�r;~�1�Eo.|�W
�W�œu[�&iیOC0>\���-���xj?l�{�r�SQ�Zܶ?z�8_��_ÙA�����zpE���C�j%�F5����+��ۯ+�S0C%�B��[szZ,e��Uɺ�����u@�������4$��^�������gzK�^+q�p�63��r}�&����m)�uq�=����9�&��S�Nk��~&M���Ǽ��_���8B�f�\C;��Ofvx��W���BF)�mP�8��s +��:���XlxV61EB     400      e0��uW�������ޜ���0s�AQX�����Л+3A��x�ݲ�]���g���#��~�`��ܠ�5������bO�$�dD�d#���� �����Ib[ݸ5��x{#LZ5��o�	�D
�@f���j_V�T�$� S�~u"g�j�%�k�K�˯������/����x���r6�VRw��,02�eSC�-}��h��>����@���j5s�	�M9V�UoXlxV61EB     400     140��jH���bE�+J�����ٍ%��a��f�_ׂ '=;����Z�)h� �Z��D���*9vUp�L������m�wGL���O���b5� L]��Ƚ{�}yd���vP�&eU����d([�$�U	S���XR:J#�4r�S�����$�3~��������#e���4I���1W�U``A�ޟ���o���F�e,#����lO�x� "����i̡���*Wz�Q���	���X��a��]��Xw�WE�.pO��W�Q"��8�ψ��W�K�N��]�c�1f$�~~�v-��Օ�
�qXlxV61EB     400     180�r,�e�r������A+�04XK�D��M��sq�|��H�Z�[��&g�[а��q�RT�����'��W�8���	�m*��U;�%��#2���/f{<��������K$*CW���9��S���BMvy��s���K���
p��c1��$�bs�[b΄:�.E���Ɣ�}2ĨU	WOJ��r���ÕQ}E�T�X�S����+����b�ꏦtgQ�Ql�Fb%Ja��"�MK���B1
ׯ;�b�36���1���;�ҐO���Uv ���Є#m�>���Z�*���~%�H!0�Q�2Ӛ���6�0;YY)�m�G?���k�6S�?�)b�z��oB߾�i`5ه�Y�5���:k�~��3UXlxV61EB     400     150k�f=�>_���-����Nv�h�a�A�T��8	c���c,��d8�;q�ʞ�z���9��Ts��z��ua�\p�5��sN����u^�ANc�2O��d��P���U;Av�}jȎ����D8��qRaBڤu����H~�c~��.8�\�G n̨q�z6
�_���y<I.����L	��9�5(�L9�҂&��)�I�e�f=� �$UK��D���8 �^XB55�gƓ�&J��4-ie
8�/ޚ��|"��B�$8�l���C �)?��7�%���hct/�Q���P'�4|h�;���y���_��֘/0�R�V���|XlxV61EB     400     130!�����bu��n�p��b�]���|T��p_�&�gW�A��Չ[��j-,<�n��^�(�R����l�xoMC��K�E�
�7��Y�X�5?i��1y�W<Y6��^۰G|��U��Ump�*�<;�p�~wRb�Ե�'���H!�Z�w��K� c��9Q�m��5�P��I�m�ncI�5�%[|�G�\Թ$o�i��"��R���{[�,�����!�.�y������y]nC�@�
��Mcz �+�ёU%���S�
�Vl�Q�*PV� ����,Z΄aVfw�b9*e�n&��Z#XlxV61EB     400     1208�<K��E�Q)�?u��|��6W�����
�n��6t�C��=E����/_���*�pt�S3aG+9���m��2���]+�R��/��tq�A��_�kީ�k?�E�N��G��:�4�sm�;���Nv�9�8�J(j#N�	'�Q��m!9h\A�s���D��^M�;��F��X`��+�f����7��<RZ�Q���cG�	�13!&`5���r0�$��q��С��$�%�7�p��f�����Ǚ[MgNiJ+s��%��je�׍*�u�r�Y1	-*-�XlxV61EB     2e8     100;W��"�ݼ�{C����6Cڤ$�W�
ۜ��8�{ɹ^�O���7�k�)�+�
}+��S5(�0dl����Q>��%.�����A�^�#\�-/G� D7�ۊ���CBpGԮ�xi)O͗�g\n��N*v��tz��M��r�)>%/�/	$�~�H@%L-��Cg�D��bxV2�\s��D��s���K
�% �y���r	ɏ7�"���G&]�/��m�Ϩ�O����/ڧL��A�+�����l<�Mu�T0g