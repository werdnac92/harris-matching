XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     150���X��3�wB�(tcH��{h��ʬ]=l)x�U�;�sxE��PRd�l7Ms(�_�S@y�GP8˅N���6ڳ�&��Tƭ�y9닅���{���],�
B�b�$�嬮!���6�i��P��-��.i��.*��s�>���6)̮g<�uˤ���x��WS�!�#KMwc�mv��k��ߙ��o��b`c,Բaf��T{�y��_��R���p���x��6MI�c7g9���I�����I�u�i�����8�
;%�B<�Cg�9A7W92�1g
��WG�Z�&�2��Eޛ��7ARN���鴕on��g9ߛ��u�XlxV61EB     400     130fj^C��W���!s�1��́6Ne�*K
j�A���&��2��I�է�ۧ.�3��E��r���\7�5��s�SȆ�T{B�x��8�,_��Edf[$?��~7�U�_����C�tv0�T����o��������q�	�9αV�h<'1jL��!��D�23��t���n"w��2��&+���GeS��xבg����urӵ�O8��w
���K�^�7�f���Mw�KwF��I�ً��t�hrH
/v6ϡ����ݯ�E>L�1�}��|��Y���WٱT�'`��g���	*1�XlxV61EB     3b0     150N���T�-��in�>�������,43*��Y+_80�O���o� ���K��DZ)s�Jk�6Q��Kiח��8X��ދ�����I�D�3�Ȣ�M4HP�!/��-�(��B� 3�f�_|u�@H40�lH�Q�^_-/��zW�|@����%˘�f��R�C̪����@�7R{~tTFa���"���huZ���ik�Y�5b� �`@��H��dS߈�\)���f��E&�+p���4�x��vw"�yۅ�e% �ꃏTohNz#Ĝ���j`��T_L�@Խ͞�=����A�ne�$8�{1 ���)(*�5{��P>��XGS���\c#���