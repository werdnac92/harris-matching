XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     150�L�¦-'B��*�p4K�)�)��VHTM')�%��ߏa�e�#�w�*}�2g�e^�rQXR���^����S��3hw��N�ѱap��M|@�Bn���5���_7�6qߢ��X���cˢڪ\�k_;�L/�֤#IX,Q;b��ϥ�l��j��s��g98�Īǚ�*�W�2��@c¨�O��ϸh��q�h�Qi]N��;)X�i?��c�'g��2�u&�P�f�~ܩ�8᷌g�ދ
�������=8��鉼F��>[�)����ch ��ɾԈ�XS�썾�`wU���b�I�\�����=%�@�Z�D���͑�XlxV61EB     400     160���4�,sO��P�#���Ʒ�q���b�ز�P��b�i�u◮�����3@�b���紉ob� �'�,a�_��/��7Ufu�OA��u��0^�"�z���@c��{��l^��ze3�3J�K�l��]c��#�R��R�A?�)�����͓���,�,Tt(��"6����0�����~ȯ���=��m�68�n�.��YiF���[��#�FaMT0{ar��o�s����7�/t�LD]�d�	ɵo��كy��8L���B]�,g�pr(;�1y��� ��E�����>�������K{-����ҊWs�-W��;�=l��q ��R
<,�_�6[XlxV61EB     400      e0q��q���ЀcAh���U��IP���Ȅ��kү��h��Ke~�ň9�t�>�t���`Ǟ��e��j���C�k�0Q��܉)���2�'9oouw��'���ͫ�3ɶ<��0�(RƦ*��^rȱ�Y3x�|q�S���<ڑ��XtC�����N���VP�MR["��:R��p��m�"���m�_�XT�3��ߤ		\@�"E�j2���fqK{XlxV61EB     400     140�̚4ɓ��kR�.��W4�ś`8�\5݌���$��8�UE%W�{��BǰI�E����DQ�������$�ZA�\�	�|�z���c��;C1^�k畈������2��x�	Y�[��K���Nub^��X�?y}���U/�/v�mV�T�˩�h_��K�²�	�S�Z[�ϕ���H7R�b\�'}#(�����+gT���#�7�˳;-R$�s?�v�Y4�Z�0����y6L2���<_%��S���-H��{�-�8��] jl�p��@P:�s{�D۴��Tȴ߁ ��5nM��P�+��(��XlxV61EB     400     110���sǯ�c���������_w��@A�5�/�9�I�� �(EZ��X!��-b��y�q�&`��<�4�&���<}�;��P>*)��Im8��:ǇJ8!*�� fm^ޕ���㝇��ˊj*�ei+�J"���fvo��e�TG����=�)��"�5�F���<�F��K���ROԐf9M�&P8.���cC������HsN�K�~�TT�����ZU��ԉOnX�hY�2���l�"�"f�Џ���H'��l�X)��h��0�XlxV61EB     400     170�ty��dO�EC���Y1@T[�4�������	���Qg�$՛ƃ��1�T��R�d��/���8��X�w��r�d�c�J�� �&���[�T��!��G��gk�����³�
e���ݮ�jZ�W����eT]�
��G�5�>��0¾�7�K��v/�E��m-���2����s��V�6s�yɏm�� �s�l}t�����K�fO���;tT}Y56U��%`�ղ`�3R��{�Q���W�`�,��E���5�9a�jK����SV$v��,��g�z��||����	/Fms>jDl�/4隸�P��z�d׶Z��=��?������p�"�M~���3�i�Ͼ�ԇt�@[��XlxV61EB     400      f0ۘҾ�sB�5�(|��۰b���A����XEt���Ӛފ�큒o0���X���k�|u�E�tWi�"�K�ۻ1�"�-�|��_%��@�Wu�a!�3��emJ(�M�x�=���)b�����֫'n.��kB�Т��{מS�ﺽ�,��Y{��A���ύ�^X[@��m���|����`��z�Í�u{�K|^��~tP��1� �9�Q�N�&C��q)lA��XlxV61EB     400     110$ɛ�)g��(T����&�3#�'�@}�	I��;�|N8^��K���jߗT�lǲ�|�m#9��*����`n)ط`1X<�FPbC�v�xa�#����I-^ׯL��.�usio�چv��zg4�ŵ��lh�v�sE�dvP)Q�;�+��]��kO��4�V�vsO?�"Vl�Yu	a�'J��[���Ѿ��9쁥�m~)��>��3)��9�ڒs<H@�i�p���5�}tI�����U��'�}��u�H�r�H��H�h����l���>XlxV61EB     400     170�lŢ�f�=�K�
���R �W38*��)��/����L����F�s&>�.��&)Ap�?���|j��2w�~u�\g^�����D� GM��^7o�(p�9A��G�:
c�N va�*o_�.�W|�C���y��_�/��hB)�%�ZrRI�b���'J6L���x@�;��p�O��Ѧ
�"�%o�1eLz�� N��j
Y����7�uǷzȚ6o�F[��9#k|5hK�^�0M	�):�p�N}T��]@̗�}<����C=�8�C:�d
�)QMvT؅JR���V�O�D$
.~��(���p9s� Ha��_���XBBC4�̲���ۏq�
|�˳�V;E=�F�2*x�	�XlxV61EB     400     100+ ��r�a��T�ɝAz�{X�*�C٢0'rS}p{%|d]a#J�U3(�+��:3P[��$�)mo�E�+
?��9�Q�^�fu
%��iX�Px��E|_�:�>&�n���{�jԾ�����4�uH�v�M�%X����`��%���7�2O���p�g̰,�0zP*t���	�T�u};���W_yf�_�c��I+�hp�R�(�8e�
�:��]ǅ)�3���z�4y�Է�m$�:a�R5�6���{�|C��XlxV61EB     400     140��PfD���񟧬����^č�D��������5x|�'�o迓�i#�5T����@���)'�޹,���
Q��_���m�$'��)���e�%e��bΦ��#s����N���#�<���X��&_�yPa �,��>ZJ���I�F;ۭY�I�!�p�����)�*�ڔ`$�j�P��_vB��uƼ$����LM�U`�ޚ��,�4�uE�p�+ψ��~�.�yQ����*(���<Xiȣ�q��S�k�ƙ
4�*���ot��bC$�cp��#\����|�F�}�sόzQ�kZ?�Q��$� Y��SC�Atc\XlxV61EB       a      20c��V��ZW�{gd�g�q���b�$vP��L�