XlxV61EB     400     160��e6�V�oL�]���C�'&" ����pe}RZ���QϦ9��2DO��S����nI#2�.^\��V*'��QI𼍧@�����mU�/��O�#$����}�<P+NN�澋�n��#J��<�󔜆l��đ`(� ۳q5��Ʊ0��8cIH�\!�#��(��%d� �b��F��,{Bc%lC�_�Mg��>\$S_�K/�ל�w�x�׾�'շ�6R�̎�A��q�Q,���i�����������+��,f�����!S���� ��<��/W.X5�h\?���z�U����z�k%�;�K��Y��uk$�b�y�m�?�s�[�7?z�D�"*��D�XlxV61EB     400     170�b�c�+Y�w�d(��|������X�[(�dZCAC�C-l �\��{%%W�ɗ���T|+�iEP����(���p�T��
�l�(�_D4 ���y�A�#�P������-h���s�mg�����3��T�~�,�aN3�c�$gJ	���!�1��;� ��`N�8�&㟾�a��T�&���q����?��f1����m/�y8�]Q��m���y��p�$�ݹ��)�*�~���ۥ|���J�����I�	��'Ø���Zh�Ǩ�+]���O��.^��S�p��ZSS�(x��E=�٣?�P�"�Y���!���J����pn�����ɴ�
�e+�
=�d�M��i��c���Y�XlxV61EB     400     140-�����G���	� ?_M0 /�!d�RTj��bw(��:ɭ�ȩ<�
{�^s_����l�ϑQ��"oQs�L2�����3mT����}^���2z�(�[�޻�H�[-�}'Dv�Mi�Zz��[����o� �}�N�M�?��{���RE���EΌ�a9j�\�h���\����f�:�LN�whۊ�oĶ�B�K�׾�V��{��:J�J����ߦl۫��CS���	���6T�f	��n!�h���4��6�^];E��}¯�l˹���|���w��w�qdm��a_�.��$�?��q�{6q��MXlxV61EB     400     190a�)�.?�=�۳������Z�����A*^{Y�Pn�x�c��d([�ͩ6���9��c����֔��I_|�|�O"`WB�[l^�t7�e.Ӯ;�7���ލ	h�	�b��Ư$�$Ar�*��Gzإ���klԥg�oɆ��|A�P|)y��W��G�J�����f�lqh �&��,�5�~�׫_vC����u>�Iv��R�Z�io"շ# T6����Lz��V��=�nM2[�����Ի��!rj�ey��`�A�0�?��/� zmc�Hq�2���#�_"�zr2��u)i%�W�r��\�^Jז����l:�*O�K>��`�c�n��=��]�m�xT��<�1}6�ou�N���g��|3=j�U7vZ�=6�/��oձXlxV61EB      75      70,G�V�ڝ[���4�@?Z�� �O�^�H �=��9��P�O�Ͳ���0��	�S�l�_2]�!�³Z�X�a�9�_��V�=5fK���r�VH�"B�)g�