XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170TA���5�ۺ�	���=�wDaۑ6��7:N4[��B:�c2���B���r��)�b�>�7F�Ձ,`�
�"E�Cb��iT�8��[�7��%d?�J�j7��Οጒɖ�F��?���Vg�F G �vv���|\����#)�+��烏s&s�ƈ%��0�)a��>�EӬ8��{n�wS#C-��@ȣ$Y:�L7~��#¦g��ҡ�|�����f	������TL^���^i�C\���:i�YgѰ��0����a�V>k�؛�(��b�*@pb�*R��;���M���W9��:ɓ�4�=��x~�	>��ن�&��c�[)TD�ppG�W�r�/K#��8!XQ��́XlxV61EB     400     150A��������Jh�C=^<�r ��ҽ�_w� S���q(l�a����ԩ�y4���g�YJ�b��-�̯ھ>�����#��H ��WdҎ�׾=+�цP)�c+�c��{�\���&�' �'��rX;,��T�}Db��M��g�����=�ٚ-�ԫ��i$���I)�C�x�'Ě��w� N�����x�ÑD�뷜���2<�&�Q+肌��6S�"q���@�Q�x�R}�DȞv���G�I�#/�űvfn��#b�����dp�w;`QF:{4�27��fx<^!���U����=N��ͯ9���+�G�~�k��X-��XlxV61EB     400     1901C���H�g��,w���/T9��6
�c�'����6!�q��W��ď������v�O� _Q�|��js��Pu�;�9E�����a�����s���X��
\���2�E8~Ⱦ�e��*���W������i��8v+Wk�!k��v��;p�M��� ˂����^�8"�Ye����bčDW��
��r+�nˠr�#��-�{H12c��B�7Qރ����O���O���Lg <��-��Z��-	�b?g��_����E[7m<�L�	A��J7�:�_i��?��2���򊔚�Y���`]]Z^���lk^��&h�2ҕ_w���㖎'����~t��}��<�.�q1`�@�r��zZ#85�~�x��^����|D�Rq����	��XlxV61EB     400     190�{��ko�]�ǪI}�-����9�/���wz�T�Ck:��1����ұ��j�zs�n��S6������8������n?�!�6~9��DҨ��)O�P�Um[=��|ш�xcZ�Q��'����\��Z�T��
�t@�m��Z'K�G��l#�}F�
�D��U0�N�tI`۱%��Ж���|��C�O�諧��ݗ�/��&�+L���k\�Yuř�^$-�-���<�D|/�M�����Hf*M�:�r�Z�*kV�ô8��Ǵ���
H��$�}dB��z��>u�o��PLU\���d��]�˽��OLr�-�u&��Z��2�~^1}���{>��
�EMCZ ܅����`�dWx���
T� B�]�-�u�zk���t0XlxV61EB     400     120W|�P��LΣ���΍f����X�$h�V�/�M<0�?�l|>2�})�q����<������I<�C���Y^CJ<P�:���k� g͔�Ѹ�Yzb4��`�q����Y���q39"�N$*����)S����STHN�xb/%�b/W��Zl���p���u����>!��>����a���җ�E��+�^men���&:'�>�C���*�����\�,� ������*I L�ŕ�5��P��^eC<ϗ��"��Hk���P/k�2�AqBFJ�x�D���"���XlxV61EB     33a     150N���~�,�M�a�y��`�z�*�I
S����o連.���7ŏ�q�j{1�L���-&�=o����q)ZP�/�4!��~���8��W;�Q;�ԈO��z�>-NUPE�7���ʊz���T�ΔXד7���J��Չ��,�ĺ,ka�4�E/�R�53,R0y�t)��>�$4�J��2���.�J:�̼�J@� �g��Ya����s&w~�������B�7�uR{g�q�S+I��|��"�Peڊ*�[���Tq�q�S�Iɉw �#E�L�6ˉ&jL�$��e��%zK�?��f}Ԟ�؉��)����c��3�(�