XlxV61EB     400     150��M��p�
���kG	ƛ�%�n�ݴz��,ˤ��3�|1/�a Ӄamy�u�>���[]o}�b�~8���J)Mh�m�z��"Q,~���
�lt@�r��8^�$�wN7;��@z���d�QC�U����m�׊��f2L��n%�wڸ'��,��'�O'N���>U��d"1������^C����9����pM���%ŗc�>�bb$త�2�d��	Y�����G�v�̣�U*=&#e�H����u�����`����|��Ħ��o��yF��֑���[�'c,Y������-�L��(��P��η���3V�XlxV61EB     30e      e0���*��5H�O��rޠޞ�!xၛt<�[�������r�QE�p�ybټ�)����T!��w��%��
פEA�i
��O����x�;;`�3~N��j���
EA M�)����1��^�6��7�^co��\�m�*i�_�]�佪dW�5;�(�� ��݆���>��2�C0��	�����d�{ʯ�i�j�H��F��P<�VI��W'Ւ9�W�5