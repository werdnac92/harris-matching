XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     180��+�Q�у[N��:����M�f���X�� �nZ�5%�`m�sƜ�\�W���{�ɖ�5�|"�*a19�9�!K]�|�KQ25ʶ��7BTb�Ȥ�=�za�ַ�m��`�P��})?�m�*�7�^��w;e�{��%��\4I��#?5��Z����}
T����~s��4]�c/�*E�{K�9�9�G'G�V+'ϋ��fd=���No� �,*O�8��lf"N�Tڋ9�D%m=
s�B6m\�|?QV~��쇞��r�[֭�>�8#�.<Vv�cpfU���j%�J ��#�΢���g�Iu�'��*���������ߨ6,�m��$_��\�=H��e�j\��r�j�0��;�?��(6!�o��6�W����#XlxV61EB     400     100���'��U	1w�9V�q{�
�f$ �O��.
�td��s��ʛ+��b���b���$\��#.��".���5#�J�I�o�~����`��7��Sړ�`|�Fِ�_/�/��~5F�G������
 ]6<�}���v
���� D�Y2�O�ZH��Q�(�q�����@��!LѼ�6���P�� �f�̱%Ԁ�DÙĈ��s�nm�>�(�AR�����������lV������J�~�A�������2XlxV61EB     400     1b0���]��q
]�P?���lY���!yDb�!m���s:'�c�߆��T��#b7���= �؎,%�9���u*w.�ü�Fhj��,7g�vr��B�Z������݋��욹����Hu>]�1�7EU� ��_���jM��Ydk��;}��f�G��Or�h�8���x.I��I�^�@�<q8t����Eˋ`aDR�n�Co`B��Zb�mJ��L�G'Ӡˡ3c��R[X�pT�1���Ԁ���V�K�4B��P_i���J�o�a��z�Oy���qK�a����`�����l�G��>��N���ď\V_�4]�sʇh���썶����G	�>�	�����-��;���5���#�BV3����p^���f�a�Z]άFN~҄�	��`���0�qC���8Ϊ��^I1�D��XlxV61EB     400     150�5��HѱP��w3s�k���b3������0�v�����YZ��G|*7��F���kW�Ņ�Y�:.9׊<�E�u�����h�W�wk>m3�Mw�1��u��%��S<��$:e����ó��QF!����Qs�ƛ>H�ہޒgƋ�;��,λ*�TXL�*�5ͺ���`��7�T�w\����#r̒3�֟n���y@��c��7�&n��<���;do�$��:wgm�x(��D5�NC��ۑ����*�`��{����F����F�·�`͠��fI3=6��Ďt��R���5=�V�\޸��H��$��B�hֆĉ�hxhڼOSXlxV61EB     400     120�n Oݵ�aP����1^jXZ��H)ͷM��=���f��|y]��&q5*0��Ǫ��>�:��){RԜ�eRs�B�Lp\�@dh�lx
vy����$��n���m��ݘ���mh�i���>�./Q�5�}�\��?��<,�N#�8��e���s�����q�Տ��l���V�(Ee�Β_S*S$l'��~`����9?0��n��`�P�ejC��p+*��m���+�ȹ/�i��R0ʹ��?\-E�*��ۨ�̂#*D��Ѷ�P��Bmɤ0%�"�XlxV61EB     400     190��ӛo���ZW�w��^8�'��,��Л�Ծ�SX�|��.;��##SH����W|F]�H��rb�ߥ24��`(5�p����:4T$\:ޝZ��2\��i���.�i���Z������E�톥W~��dH}���9�É��7q���j~�_F�DZa���C�%�lA�4E�
��d�dt��S��_��p��br��l|�zS��Ų1ޜn�T�YJ3~/�ǿ�������o��I^�K��z�ʥ��B�hd� �gV�6{�4�I�I��0�j6�)8]ޯ_s�';�R}7G�3�午J#�;u1ɆYO���:[\}2FZ�ɦI���G6���Fq��X���C#n��I�p�:u�+�+�����<��3�U��|~�&��Q#x�-1m�����XlxV61EB     400     160 ��h>��_WT��u;q0�}{\~�GF,�/��63�N�S�v��嵐��� ���Ճ�FO̺��9S�1�卮o�[�	=�Ѷ��C��K�Fu��Bv�p��Z��?)�A��*�����w?�c�\�(����--O!-�h��УqPֳe�
U01��(3����Y?� �
xX��BIJI/i,}c�����-I�#�����h�a�5���6}ʘ`��rDp�O���y���Y�6萻�� �62��i��E��\x�e���UѠv��>�y�b��<o,4S�r���6�+�PP1�EV3��ݷ7�Pg����Pu�������|L�ȩ~o҅�e�XlxV61EB     400     190���ov��+��++�9��wR��:<��u�2��a}���0$�|PWC�ކM���NG[�xo�3q�́d�`;�`OZ���D2���S��NӃ @�C�,-^����L�e[�cvj��ή� )6�YP���+���V��nV�������[7��'��P�q�)����,gM���o�b\�(��J}�dq�ߝ�8NN��!���L���պ��|�?nu��_ P���I(ﭕ�؆�"��_5�����Ci�Ș5�>B�������T���_�a}yc�,��ޱ*tUJD�����O"�7˰ۦ�S�?ڵ�}j׼R?�	HHxH�.�5�'�|�r���o�����̽!�SR��D�6Q��s[#�q�#��y������	*�	{E��}XlxV61EB     400     110�؈Bk�ZKG����l62�rǒ}���Q"{���u��@�i��M
��z�
��8�'c�uZ�8�4��M,nH!����nxn�ǝ�"ly������y���)q�(�F�WC��0�\0S裝�!턐`3B1�'q����!����3�ߝ7���+/K�!g��nZ(Sk䣂Z-�	3��X~�ܢ��5�IL�Й�-7�-v�d�ng�Q��P�<a��0U=�j�@�B�3d���
��Ae���76��BT��?��x�,*x�TA����XlxV61EB     400     1904r��XA�?L�NڽM�EY����k[�L���mþ��By-_��'=��N@P^���_��Ҿ��`Æ�m��`�a!sa��PL{fE����A�!^._�x3W�ѿ���������)'x��9��	�Bi�1��߷W�cU��F�Q��>q��pu~�MW�7*����ʥ�Y����z��AWy�i��N'���ߡ|M��=�_��aT�S'�@ |T�~��T�����n�,Dl�bJ0�xjB#��~��+ހ��c������>M�G��5����=� �z�qA��DE�B��ac���@���/<qy�	������� �*�H�e�XjS�Is��D%N�-����?�[՘x�q)KX)~@�!\�~�pw��C_eżZ���!f��XlxV61EB     400     1d0�&��j����W�&d���H8|��S`>�����}م}�����\;lS��>%��!�ߚtO�j��p�ӗ�5�18m��G<.�=5�kn��O����ꃴ
@`"y��u�A8n��7�,�BNpD�����y�9)S���q�aJRDb��*Z���T�� �74�Gn�/΄��ڻQ]��uV��*zT���V�`��� V�e�̟@q��m�0��{�1��~ʁ�5��ݵ�X���e�߸�4�fgp�槮�Ԙjy���Y3�1��AħP�	$7\���|��j�� H����d���R.�W��fa�X�������hПԕ�_,�_F_���Y�I��;yL�5�c�N yQ��:��Yg�6h7~����EM���J��VYm�($ϯr���D���}oQK�R�y���[L�h���-N�Bl���"���w�8}�`AGl�wX�����c�J���2�؏�XlxV61EB     1e4      f0��G�&�I�lP��b+�$�x�ɔ�e���.��,����	_�r��2�[B�\�>	s��ļ���)��n�ZC�~Li�r��_�s�d�~u�N҇z�լ��ȷ��F�`'�1
����"�{r-1��T���jf@�i��۴���=�+ ���h �K^����5�T�ʉ���I���&=�u��O�F�߳�w�C��Z�<��s#�\maW޽䏪�*����2h�X