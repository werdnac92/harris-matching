XlxV61EB     400     130D9ɛ���l�k���G�b3�sq��$,�:�� ��n*ٖ�R*�Y^���8��S�C�ME���k�e��H�S�5Z�F7�n�0�nW�g='��@�vL�e�nm%����`�a�'n�E���h��T[�v��/U��#�߀�ǆ�^���e�=r�3�8�5�N3�2h�
?Sx�w,}�?�\�^����п}y�%8E�d��@��=�g���րO�+V�0����=��S���4�;�յU�o� x�'VЪ>nS�*A2�?�����fz����p�$eN?�+屈�ߔ�(WXlxV61EB     400     1304�[U�~�e�n�Ո�N��oLSj�i�St�h[��=8 �}S��S��G�n��~�:\�r�}7Nh-�	��'������(�㱞�U�ʉM��&�qy���v�'���׽�&B��������'�"���i�����=)q���{O��
��V�yBTBΛI��h���7���*��}!9��h���� �K�L���,�MJ$є��cY$Jq��Ǻr�E7��I�tx�F�eN[�kdH��W�u�1�YCfǾ��#��N%��N�Q=��]��k��ȅ9�����H��1XlxV61EB     400      d0�/������$�")jao߿�lg�%�K$��"�П���C�}� ���k@x䇮b)�yi�<��N��5)(�]�(J��w��ݽ�5���-�xއ��E���sk*\��>��2kSΓ��*Ѐ��}��Hζ��J�t9���=�`�Z�<�J�/ڕE#�Ƽ�\x\�±G��2S�c�o��92M"�,�Y�XlxV61EB     400      40��<Ɖ�����H~�` G�f�=�(�\���i+R�!,���i�N�I/"�N��$�X�"��"��XlxV61EB     400      70Ap-eb#`iR�g*��|�$���<h��v�����Э2ǆ��� �3/��0�;�W��Z�&I�)��Nh��lw�/�zG�%_b5�7ҥ���쬿��)�j�M��XlxV61EB     400      80����~����:V����uLJ����>у����I��g���mX̱j���UX�^_p�R�6����<�{�zQdLء>�G{�Q�	%ׂ��Sh�\�_���[��"w{��k��M$����pXlxV61EB     400      70޼��P���{>�b��<^�	��{gc��zH��|n��q�8�uښj7�y%V�s�#/�(�H���g��J_ ��U|ɓ�����*��T���D�NO�J�WQ��U'�O4Po�yXlxV61EB     400      80�oF�1��=�wH��@Έƨ��曛�K�F�it�w�2�}��A��5T��?�q����_A�F?�Ȗ_��!�#��ꔬ�j�� �W��b`LyRRﺌ4=eL������Z�ˈ�s�/�����[�XlxV61EB     400      30��l_��gr˸���TUH{���{�P�ݚ�ӭ�F B!��}#��?XlxV61EB     400      30���;�~z�%z�u�
, �k�G��s�`�o�h� ���k�x�!�XlxV61EB     400      a0UKp���v m��x����v��)��U��8=x/w*|r#��5"Nv���jĴ�~;�I,f{7.Ab����_#\��K�-W������i���r�/>�ׂW�����ZU��E�͉����>�@ۄ�ހ�M�sB�">���>ܿp�d�n�oF�$B`gXlxV61EB     400      70͓ޛf1P7Ɗ�0Rdm�J� s?��*^S�qS|����1���+��¶Pt�{�RY*A�7�$��|����� 	$��<�A� H������������V=��L��%XlxV61EB     400      20�r����`h���7�8�ґ���fG�Y��VXlxV61EB     400      20���mT�@�v�#�h�mO��vi����V�XlxV61EB     400      20k�|�Q��53�9Ӵ��e�|�8�JI�d�R�q� XlxV61EB     400      208䓜���M���۴[n�k&)%��¬CJb:�XlxV61EB     400      20-����*r�l�t��잲�	����dM��[OXlxV61EB     400      20*g�N�� \d�3vL�
S ����-1l!��XlxV61EB     400      20�Nl��s~['��:O�����w *���hF���XlxV61EB     400     150���d���꥗�P�E#�Q	�����}�5�~����J!^�W����J��yIF��)�x��+7��3���Ř@�>��S����U9�تSE�Bq�ho�=JW�?_PT�(��;|vN��ن�J	b}�Ӎ_~�u^o����1Ȫ��\ �٘��ъ&�S�����n!h_�M�<��;��8l7sL��Uq
5�6����=��[�k0�,���3�N��s��_Ȑ��JY�J/�/��T��^`m�`]��T ��<_��"��G&N�a��=����g8�{�����Q����{
ur䵵�S*�[��q��e�S�_��!H���D��XlxV61EB     400     120�����w�a���!Vh���(�l�6��+=t,h���GDk��1e��f ���0���ɑl�/"���wW�N��p�[ȣ�]����!6����h���i������Kg��:jb֫�-N,�^8�ĵ��ށ�6w"��w�{�F����H���]�C̍{46U��kHm ��gS�L��eD'ͻR������G�`����)�<hp��0��Zg��Z����%5�Ә�*0������E1��U�. �_�R�<h�U�&��Zd����9��E|��,{���XlxV61EB     400     150��Y�V���#�r����x2&��������{-�T�_���]i��1�S�Q,Qc�8��y�#Q ;
���؏;`�:�$�Pr
I>�x���=Z@n����^��mWv	�A��/Cv�S��6�XI�,X���ל���&��*RsI��,�o�('�}��5�+-�h�_^�u)�-'���u Ȟ	ͣ��}�9�i�L0k����W&��09�,T�<�+�aLy�t��.w,�(,TC�76݂�m"�Ǧ��'��2�wc�ѧ(h�Z�RL�)��*[m1(��ˆ���@�y�o� �\��[��)��,;��A;��t[��)0��{9uXlxV61EB     400     100�J71�#v2���w�F�P�$��Dj���1�ۘB���12�(����ά�6&r� L2�ޜK�-�e:-�@ܹ&x�k��/��,"fWo��{�D�+K���<8���^��7�|A�M��T�G�9A�6��?�(�%;#x�޵.}����Dz����c�~�O�:��]"�yR�����0vB��	��'a�<~��S�*����f@$�@4�Ou>.ѿ��n#%�̍�'dS��z���a+��K�����������XlxV61EB     400     150ˁ\�+��U��NA�"�
\
,,6�vl� $;��zW�9��R�t��;ا��TUZ��^�X*�
�į푹0�ſ�+�LɎ�k|��Ta�>i��G���{$�(+�k�X˒s��Q�4�g��*�3�����U����J�}l���4"�#Y�F	1E���+���VC���]�'����i̜|~ÀG����0��<'z��ē�o���V�%�ٓE
�
ؤs��Ͼʿڄ˩�A'��O��y�?�K˻+���O�N�o��î�e���ΊبOFEθr1���M�ų��.�o������i�=;M{�����~	k���&.fH���TXlxV61EB     400     1a0:0x`#��%�~3?Fa��K������<e�OL�ݶ,��$}�/nY�i����հ���Z.x6^��h��7�`�����H���1�`H�r�Y>�����H(=u�~�#�G3ý��l�J����p)h����
�\�ڼf>o�؃�$B��s#q�ɇ���J��K��6Q� ��ꝶ�W�@- u�1&����['�M6db��L��jS���[ϼ�i�/��-�:P�c���U��<Z`��<&�c��%�u�W�P�8��mWC���h�8��j�l�i��(ɱ�8/J�V\�	�d�`~��f�pf��u �}f2�+Y7D+H J",~�޴LD��5�M��*�+T2��=����6�oC��=Z�TWw��K��hX]#�V�J���C���!"A�\�XlxV61EB     400     190�@̂�V�	�]Lj���[��z9%��l+�ɿ�H�"ؔ�hym�^
g:/���o�=���^\G��a�~	��3j=���e'׹��������vD�|�c�����p�h��v��y��}]G�,�[l�tٜ��x�ZO��xQ �H��'��2l��ۛFA�>�5r��hj�9\�ONy���(�;-����_S�1Ho��8 ϭC�\�k׃�XEFD;�hR���Y����Lh�/�֙.��O���ڿ������t\L'o�ed���}W՗Qy��7�Fȋ�&������"uk5�%E��L�DjJ����6�
_H�õcY*�8�R�D�9S��ш�{g�JD	����ss[]M�P��0�aX������Xu�^��Y$���/yXlxV61EB     400     170��xB[��ҧL�M-,7i���>���ܩ1Z9!��NN}��o��ŁsG��f�R>J�7~��|���$0�a_�����_$����V�H]�s-��郅/���._�R|j�@��q(��{�	��ϻ�̉�S7�Qe՛��&�ay̩�@Pd���ii�������,A��%$#�R9��ׂ�X����T�k$��R��R�>�/��1w�ߕ�w���T����Nd�
J�X��2�񛙻ʫ�&Ecgx�>��:�-�۶�+�>���qB�րk�8��}]E�@�	;�V��#Q�}��i�j��'������� �i�:Q�l]�3���1���[��Z5	�6ߢqxZݙ�j���DS��XlxV61EB     400     110�� ��Bi9�����,s� �%�F�nC�<I����YS��f%�zcR�JK�!���fMY�,.rs�x�s�}��yX�*�rk�U����k�����g�xP��	�
�s̼��e����ސ���^���Pe]:�L�[�Ì�ё�z"�P��X
�J����P��x�`�j�(l��\v�_�m7�� tܕA�>,�z�eT�̺���� ��\3,<�ߧ2��`9C�~���ԏ�?��蜈(�?1!�:���$�Vy'�aY?ӈ4]���XlxV61EB     400     110"�u9�0"I�� H@�r"�@�2�(��
�X¹�Ne-b�.�Z®�y]�g �X�����ak?Kq���
U��G/o�\gr��,�H�2El�@ڥe��A�b�5�W��'��7��u�N���A���'s�Y%S6�	����o�z��D�9Z�1\�;��*X���MLVL�Y�����Pa/����0î���%b���
pV��1�⒇�RSG� ����ӓ�{͢B�;�u��:8jmI���L��/���.vn$a�|�XlxV61EB     400     150�T�&��]�1>��.�Q��͝���;P ������u�n.�]G(DLj�PV��3h�����Wr���HLS���z��v^�׵)���)�Ahu�4���F�D�bR��<�gƚ�����'�FA[W�d�g̭�2`uہ�K��xo�*�ơ�¬�FJ��-�oO�ꮆ� "ɴkzخ���ǔ��SiG� �_G��8��޷F�G�� ��I�M��i��Np�Í����]�g��1A������a=��k��l�]M1o�^Q�=/�||�U2�'5C��5�����|)� �;G�d�������'Ǒ�A�XlxV61EB     400      d0�c�K柃Yw�2ÎIW�k2�~/s ?�	�C��\����Ѹ`�t*M�Ʋ�
����,�Pe��y�Â<�ɳ�����?���D�H-�j��g�
&�?q�H^R�H����t����"%L�s�	�*�-�����g��`��q�����`L_U�2�Xfp9��xB���+{Ea@, �!�+(V9}�XlxV61EB     400      f0�e"ЌN��7H�^FɈw�[�aӧk���6L��ն�|�����\�T�r*#g[��RJ&r�����'�	u��Bn���:�K��G1(����p�#���د]"���#�|����Iw)���X��5¯|�&C	��C|Z&����\���6�j!C.�@�P�q�0l[���?\�!+[xf�������ޏ븶����{f>��sw�t�y!&��`}�c״��5��XlxV61EB     400      e0������p�"�\���T�<���|'J(G��L�+�<Ã؜J�Y���w��;N����yU�Ũ�!<~V���7?��=����qn#��X+��[p�%�ꐭk�>�8Vݷ+����E��p���('��*��2]�>%��2J��:`x�QLܖ�2�ԏ�0+�p��;�|�%컿T�f�*�G��y��Q���L��ԩCڥ4F�_7XlxV61EB     400      e0�=��6��(�E��� �/�SWDnD_��}n쮱�qjE�9KB)�*��%v��lgs ���$�/�/��h������*!�x����X%D`����m33U�MD�����A����|iB�1��P�m+���j{��2��\�����|aeٞ���A2�{Kp��֢�h���vz���Z�=���@�Xw�ڨ�7g�H� �W��������&�u�؊�����XlxV61EB     400     130�#�>l=۴�m#��=�"c�e��~ONOqD����ZlĄ6�9B5X�G���l��ݏZ����'�rί%�{k����8��>�x!a�ׁ�H���%�yF�O�`�L��-{~:��^��R���#$-����)�ŷCD���'�|�����c?q��m�O^gs�!�~uZi/]UJ<:�[��f8�U�e��Mό�W���қ�Sa��@K($���z�D��k���_��ט'}A=~�~�NS�
�� ��1\!��']{�y灾�Q�Y��0V��܃�x/�V�%T�f�m������XlxV61EB     400      f0�X{�;Q���Y	X���K����i�sF~|!fɔ�f�~J6����wI�ƌ&3.^���b�x��fur;l�r�����y���#9�W��$�ᢻǲ@t�"k�;C�^!-�F{�%�=�I�HH����7�0�1��5�g����Ϊ%<�=F�D/��u}�RvH'�C@v�KA���P��� ��\�s��F���ɂi�M��}8��L-��ByKiv�o*#��}�1��XlxV61EB     400     110vW�-��{39��So�%=(�G�_1���Z�I۾����$tng#1��*���R�,�!�ڱ&(�X�v(�2�'�}�G�����@��fvRB�k.��dЯPiwH�^̫�W��7L� B-R+Ή�n�oyN��>��*eX�4�P\�=��4Y��h!R<f~}h^"�+�s��9�8��?8VzG�k�pi�z"�S|^=y�]h2<�_1By��E_��_'�K���s�����_0{� ��D����$,�)��M�E�UXlxV61EB     400     150�c\5�P��^�x��7/�D!�Ȉ������(a��\�l�����k#�[��nx����Ó+
�뺰���N�#y�Uϔ�DYhA�B�]�E��g��^����KP��C�.kh��4|nE�<&�؊>�=K{�/��P&�y���Jd��E�H�U ]�<c��	i�xC��I��w6���2���Ⱦ�Z`��4Ƚ��P���V�GC����,�s������z)��$�@�������C�ܙ�)[ VF���j���߀<gJD|cF���5�[�Φ�����&��w����ߋ�Ӂ����"��Q�J�`��/�3?iL0�/�r�m��J>R���XlxV61EB     400     140�5���t����eOw�pJ���6�5ޘn�h���'�D�����"
kԺǞ����'�]������ �4Ǜ⤯ȷ��C��GT2D���b�dH�C���F���Ã�k��X���a� #g\N�ޙ��%:�	�EH��R������+D$E*�]~6}L�hS�����}m�lJ=�nm��:�7
(d{�l�D��ڊF���$�O�)1�
#}�x�E�� ȺG���4��*)��7~� �A �C�Z�_�#x֦&��uI�R�@*f])j��vW¼N��u_�oy���C���������"�'�%�{XlxV61EB     400     1a0B����N3�`/@CCx·� Y;�7yuc�1 �%��r�-�Q9�S8<�\���h�� �mvO���&�����d��!�ÇV��Khgt���$E%<͝�y灵���է�㽞c�h1��d\�T�ܥ�'��x��vɭ��=��/��NR])�d���m���$�W���j�n0�ᵫ�3��WFk���d�K7�d^��;�z���v!���q�H|�a��6cM�ߗh*��ח�9�{��&�z߯8��g��6߃���I��+����r�8g�v�`@�T����O�!^?���M�r����Л��ʯ(4����(O�Gi
���/D��&?'�a��`�;��Wk�9�������ȦՎ�ϭ�o�l��"����}o#yS�5\_m)2u:����d�20���I�XlxV61EB     400     130I��"9x����̣;Zf��7��w'�K�gU60LmBי<F��H�
���t��Q���`)��=��1�c�('���t��2c8x���&����1&�X�*r&_�����s[�H7��S�YՉ�v�-l-���g�O������ ��
�!G�����_���"�h��aM�����4��V/1��Q�R�L�xؕn��O�[+�N��nh���v�,d��[x�g��y�SI~�Kycn�lJi��&Fk�܂s7xj���<��%���]W��ͣ�<���`�}���I�^�]ؾ2�Ċ��XlxV61EB     400     110d^��reqeM�:f�\���CBPL��H�w����OnG�%����>�j�1�:�/��ƨKA���tLDﴬ$kt+���&^��,�~0����V���qx`cK����pG��#z�L��H��F+oI��T�?����6ը��1���~n ���I�����
�{��yxNr�-�hK／��1+���@F��%�|ʯ�%�1�aO]�s2Ù����QX���Fo:�]�&X�,1�L�z+̥�鵔afݲo���I�zXlxV61EB     400     120غyO+��4C�S���\���p(�X��T�>�Q��!�佺�fO1��:%��(ڕKA�af'������2�~m�<G��{��l��fZ\}��n�������c�⿨��%wc��)�@JW��o:�N*Cc%Y����J+��S�"�}����c�\�&!O2)�붕4{?�����+�����U�G6G?/W6%�ȴ����:�2b����\���X�H�
}������)��T �g�3�{?�7���f@B�D��	��0�X�z/A��\�@�XlxV61EB     400     160�,-O;;��.���T����o�A
KvWH��ow����@"kO/��d,���S2��a@!��2�bt�_�荺m@5}��✚~ s�e������GA�5o�C�l��f�{�6�r '$���JZv�nF��[��7�Z�0z�Gjo¦	#����n@Q�ӝ/��.]<��Q��k=8 �?@ʔ��7�zP?f7[}�{�P ����ǫ흋�B~Z.�r�eo�d�6L�k�	=���Ќz#/0��+c�نR�t;����%�uN��L�p�*�o�I����;�X=�훹�\'��u����ޯ�u��D��p�n�yؕ$�S<w��"kwY�J�f��jy4�XlxV61EB     400     140�%9�l�l�	�٭�;v+@y�F=�H��Ey�=FȢ �]ӢC�G��~��ޔ�CZ���F`�=x��J/���|n����a�����3�B�w��� �eH	��G�?�8�RS`v�\q0>]𜮒�10�&�G���I7�A����@6If�����尽K���M��ߔ���ݼ�eL\\A��h�3@{���EJM,7#%=�TONh��.ƶ!�g^���5���!Ri��Ibz�M���eW��J��Z��H�8����0y�m�5e�7!S:uPTeu%
��ľ_��;����oҶ9��$l̮��ռc���"يXlxV61EB       e      20l����55R��rh���9��!H�//42ZE�uw