XlxV61EB     400     130��M��p�
���kG	ƛc�r��j�p�YO;���AĜ�/���%|J��YH/]R��i�y���7�R�PrЪ)'�̬N��*w+���8����nVo$N��:Z�h�S^<�hg,"�b����7{�;�3p���lo ԋ�"�/���?�aA����+�����~��K}v��00e��Hw,,ک����.x�P�����*�;"�Հ>���	h�G��� �5�0F���CaG�E����XG&�����m��bΝ����X:t8s��k��z���G�p��Ձ7��AW���XlxV61EB     400     150�3���9O���|�����Sh�=>J_H�/%�Nt*�$�BZ��$$��G�q�9�ͮ��>�/uL��s�����$<U�`퍈c�o���Y��#�I��g�pSY�zUn�@�p~���2y�π\c�=C� ���U�V�|O31��V�u�F�qY���3�$T0d�J'VY�:��ԑ2X��~����ګs����|K��4����C�(�38�=�T�\�J76 |ı��630Y�p"���c���T�u���G�k�tA��^S/|fTK�c��"����?n�� ���a�B�H�H�vw?̍{1�2� X
��{Թ�XlxV61EB     400     160�_����"��:'O�Ke�x�gQ0�� {`M�+^iv3��>B�b��gť@�gm���]��ƒ��^�W��;/�v�W�E>w��5"�/2_\���;n����e"9�	��e6��kxR w�,h��t����Hz�P�{B���y�5��j7���q%����h�9&�r�D��`�4 ��ڸ�^?{?���I�D���9 ���^�36P�C�b|b1��C�XR�#=�v�KrX��|&y��&c������מX��YvRۮ�s��JH�����BR�0��<�c����@)�4�̪�2.�+�
嵓Hz)R� %���3$��.&H�E gW�6��XlxV61EB     400     100#vn%��:޳ag^.�)u��Je:�D�U%���U�N��Е�e����B�y$�h��e3�r�
f�Q���^JFV�h�Ev��E �)~f�P�:h��Q����ڸ[m(��)��_�zw/�P�"��43�`=�8��5�U�yi0����˹�?�Gr]��A�oSC٬&$�s��^%���Lq�j�Ii������.�B�WA+�J�=�ى �Sc~Ⱦ�����g�>�J$W�F6a�LԐ�	�蘉j&ĴDkU�@XlxV61EB     400      d06�x�)ؘ�W���](I~��%@��n/x`I n3���9lגA�nmǒ�6��-��OԶ���Gr���^�u�=��?^����8[M�o�^R���k�eђ�����"�}`���?��4l��q�,�༟�S5*��=b�S㋨��dS~�h@�qU�}�1|�F��׈�QZu�uB�'�V�w��ӕ��Rl���6Vw�2XlxV61EB     400     1600
��.�����N��ǭ1_ּ߲JM�\�3JuY���M'!���2 �A�cT�V��0?�e��[J�J�__��1�m}����?�+)��c�ե`�=QR�_}�}<du����n�\R�v�W��mȂt/?ꗿ;�x�悸x\/ze����G����%�YR��	���J�Do�)B�Eq+�-=p0]��_��7J�4���9�nt׼F21(�Q����ԤL��z�l�
~Euv4o��ݼPFO����p#h����
X:EՔA"g7�6�����/�h���'�	�J���a����ʯ3*�����w���$�Yz�-�����E�V��ܿQ���4�!���XlxV61EB     400     190�W\w�sAݑ��<�����!�Ó�B�w�(඿E6�q�z��&���dQ�?&	�(}s>-^p�!��Vpjqi3G�2��IAB��=7�vLiӖ�*�[��,V��o�q�g9U��@CH�/M�p�?m,�G�c�Ù�S3ϐ�G0�ŏl���=҇N|M �Ԓ�r�ފ�1�G�S�;E!��n�G��慎�� �FE-�S��j�/��~'�p�;[n(�
���E�}�U?b2��d���P�Y����J�ʜ�!!QE���*����X��F���L&?�b˓�$�+��7�BW�;߆����vE������=�B98c�o��/��@�7�����}�D���LqK�A�����%1F��T�f$��{�W�<�
��tXlxV61EB     400     170sK��b8���>�uF�4��R�"�!@N��uqQ[��V�]_ARl�a��/�+]��z��Y�d�ϧ�&��,W}�F}�;�6nG�P��Ο�&PB�i>�Ϛ�k���Ff��n�]�����\����Ø�����Ɵ��J��Sq���� ���6�md8��[��h����!��N�����)�/ۉ�~�.ɗ}�F?w�0��:2O����K7_P��2��v%�!��^��B���s�w�)����E1����-lEŗ������d�<�6)�z��O�ў��6�1
w��a�%��q V���q^�鵨���w��`�&�a?O����A�m���[���~M�AH&EXlxV61EB     400     160��J.�+����1���enizG���B�,)������w�?�ʁJPSH"n�3���3<��M��D�2&,̍�,��L�@w��?�Z��^�����j��8t�a�.�����'��_q�X�E�k�L0�`J*��CJȨ	���E({
�&�����i���� K��	�	����{s� ��58��m��7�	6b^�@ŧu�}S(z��N��["�����X�Kت#��E�J"�Ot��NI���\@w;I��xa$Ǒ55�ӽ��6f������K;�}� gŻJ赧�Z��&�Ь`J&ZCEh#��"�uH[@���s��8t#�Z{a�j����V�m�%8���:�k�URM�j)XlxV61EB     400     150�VlZ?a�iy,�uHL{Z��?$q�to�~���X@^g
�.?%�aB*:i�|[�׋��a)tU5ƻ�{^]D�ۑB����: \pu���0P'�H���`�W>�P\䥀��(�IEj?�pM�	��Y����tEx�9�����8O���w�"諟?E�_G�σ��t�^OAi9�\�5]�%�S��xV ��[�Kbu ��0�=����|� 
 ����M��EB�M�����^���}g�*rމ��ZkÀ�ܼ�s��;z6��J��"��}a}9�A&$��0�:��%!�DeN��]�F冺�k���ݯ�e ��2[���u~ax&/ӥ,U
�XlxV61EB     400     170�B���U���FX��]>���z�Y��d�	]�^^X�/�]�w�yӲ;:�$�?���4��jc(�#�W�S�~��O:wM#���A�N���!_�4�r���kŤ�LW��ɧ��Q�0/GA=ʂN�����9�?m'b)Fމ�daû-_�G	iM1��;t�о���2b�_����{��h��Dd#z���t����`�^ZL/u!�'k���SKV�O���C�,R�/�r����!i�����c�>���fd.�����qY?�V� ӧ;��YS��I6���XW�ߔ�aG��X�7�~5������1,�I����-z�8_2�u�2����<e$q�if�Z�#�'��,9{ ��5��ٗXlxV61EB     400     140�U����r�az v.��5��S�4#�(h�R��e�aKv\�#����]�V��Z�S����O��O�pH�Ch�$����a��B`�`�e�ݡ���Z���g`M�!��Ҋ��®*��ӡ����F�x�b�Ф�J���t��
I�2@a�ISB�V嘮G�8T(!W��v�U�.��('M��s��#	ba��+	�u勄*��49�~�wCNb��֠Ek$� ��IB�j���ƽo��u��}y�jh-F�?����#y�[,���X��9YG�U�ר����h��.��g�ӛ-��=횐�
u�v�96���B�Vs�r���XlxV61EB     2ba     100f�#P�as�'�Y��022Ĉ9ݥ%�1,�-��P�S]m�Ѽٖ�.�� d(��,�O�?�-���d��4q�'K�7�.}p��i�ӹ��&H$['�A�����
)\wIA�6M3�c��K"�^t��}&8�`$2�i{�HCa�w��>td�*,�Ϸ��0`����φ�o��W�2���:[��bo2�V#Z�p?-m�/ �:;$fJ����z>��J�{G���뺐��� ��@1N=�x���y1͋��