XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     150��kC� 1uBC��Cn��a�M��H����~Ŏ�����HӲmѤ�k��������f������IT�����9y��m����n�:�?�vm�g;͂�+M|�K��57�Ъ�U~���?�ݷ�P�/�^��`U{!�1;ƴ�=���&��B0|B=��m)�."�G����m����v�>��X�_!A��?�7��C8 ����N.���҃��8A�!Nk������Rg���q��/�zmp,�ֆ�qQ�rhK "ʩQH��}0��m�O��]xy�ГM������au�;ɂ/����]��<Fj��E����&+�/�.,G��Ӎ�VXlxV61EB     400     160�t�7<X?���Ik�솸&�o/�x��p/����x}���}�84XG� �J(��ݧ���C�!�ԬU��6v�!8\�]l�'wPPF�0I#�/�L*|`dsEttd�+�x��b��+/�C������Q�w�kUwH���Ķ5Y3o��n����jW$ͧ�X�J� �F���;Ƈ��a(���>\��ZWeC�~��!b+Q<آ2���:*��f�	�[�$>n���i낭�	�Gl��.�I����a����	V[���ӯx t��q�n����N�IK"N��?��W4��d.�$���>�:�_P��d����+U�9��Ȏ�ξS!����p���XlxV61EB     400     120Y"�;�PCuٺM�,���f3�VR��P�s֩"�2�*�t���*����ׯ�R{��L�٨�:���t"kHP�?},bw�\��r��:乩ͮ����P| ���/����̬��u�� o|ԗ ;zIo��^B�/���n�{�?}d����-u�^y���������{��M�{#��$F�P�_K�����0�CG=E.�����ȭ�َ��1���i�>"o-{ j6�ctI�+�E?��Q�!�����Nn�<�WE43&�I�H� !NjH�E�ˎXlxV61EB     400     130���.0]G��O�#=m��ĳ��`(��]���ޭ�h,��©����Qh화䵾���`#��Z��>�0@b�Q��0�ojhi��З�p�[M.��YNJ�V�Jv��@�����0Ƒ����~�W7�eZ�{m����~��X�+��^UY����=x>{�l`�	�cp���
H�v9�J^�o�aio�������4���Tv W~_�P������������<�嗰.����������G� ڳ�^�>��6'ʹ$h��V�� C��K���[�������c�ܸY�@�ܣOO�U>�XlxV61EB      de      80r�WW���B�����@_��%^�-�,F�0������t�pi�p@��ĒN�ۻ����g{\��P4 U+)�.�aO���H65�8=/f���/�p��Mc�-�f�l\�(���O�xR�