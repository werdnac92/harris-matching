XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     190wZ����Io�Ʀ�����*'P-e�T��d�}΅��������!6�Q�$�k�"�\�-�ª��1�}#���D�����-JJ�}$Q���� ts`�m��mH/ٰG0~���x�X�(�w��
�J׻"j���Y@��A���]! _�����cP.���N��I���w���V�,��>����Dv���z\�aEj&  �&�E���c�8�&�Kj~��;���'�0�W���ͤ\(d2&���������@)�Ks��`���M�I"fJ*^U��+z�\��5x��̩���������:n�km�ۍϒ7�ˑ�W2���)@�k#J�$���`��d"Ի�?�	4�=I�=��_�P^�m0�6M�cj���i��_ν��Y'6դ�E}�z��>S�]��XlxV61EB     400     1d0'�s�|�D��\*����&M�x�&�<a[b�
]�/%�#��l(+�������s�(�p�<�����X?xk��=,�k�ǽ���&����*8'e�-�ȑnbD�����ڪg.g��/��U��_3�]��\*E�i��Q�~cx0~_@�4���'\��.���#����i��He!���UVN����<�V���&(��;�0�1o���N�k���q;����iYϿ�56�=�6��W���[�䎭����n�^]�W*�g\�uL㝄1y�c/�C�C �:|�!c@G���@q��r�O�;�&k�"�vc:v4��3t'�I�u)�P�x��35b�$�2�m;X��BCϝ��Oɉ��G~�x���F(I���e�]#%[�[���M� &��q�Ь���w���2��؜�J�e���/��D=��<�н�XlxV61EB     330     170ׁ{�z��c����s�4	F���l�壬��v�d2�|��^I��8��Sq�;��Jo�S\���׷�g���Q��������� #�7���2�+t�G;�^�o�bs�,[>ق65�j�Z�}-|�JBϹ�q/a�s�8H,E�`/�L�N06v��GYB�Gu]Yq�*�$�7=��X���Z�?l�	��~�K��e�FL���Z��;ܺ�����)�HY��PWZ}zK��*=�2��?��g[�@�>8}�]l����
�Ik�Vy������l}M�;i�p������F��2m��g<�s�cݳ�e"��ۏ^3�{&M����ߊ��#Kn�Jd���Q��:���