XlxV61EB     400     130N���1���b���;B�j�#ǨkX��;qt�^wɹ����7?�^��D��x2�b�kB���[�����~JY�i�B���Ou��dS+JIE�9�,��R ��S~��}�`�34#k��0�و��*=e�J��߄Z�{R�O)n4��]pC{�����4ୈ0��h�����y�*r)��<!՝Rz��[q�@���H�t�4���˙_�"bN~�2ƓKM����\7F�$a�uM�-�J%iv?�ɔ�	���)���89EE��D-�4 \A#mS_�^]J��Uj�k����XlxV61EB     400     170�Ri�R�~��ZT1wPt?լ�N��Q*7�t[h��2�A닠�� z��j�x��D,Ĳ�>[�3Hej�������z��Y�d�{&��-]p��_�M*����b�I9]��d��;�@����R@�(�'/��{��8Q�(:r�^�~mԃ@WCO�9Y�7�����4��0W0�MK|v@�E�6U�`��Af�_�Z�� 7��^N"���G�����R8-�Ԑ����5����6����i����Z�y$�G�����d����:�{ჯy��r�5=�	8o;l���Z�w,?/���!p�cƄ�oM� �"f�d��bˈ�O�G r�������r����ש���:2�b��c$O)XlxV61EB     400     110�܃n��F���FF��\('��cN8�9J���"Ґ�ج��rI�hlx�ٳ/z�Ђ%F��J�k��X�R��.`����lU��R�dQ��͠�b�KQ�����I�����	�qd'��5I�v@�?Vu;Z9�1Ȓ���5�8�5M��:D����͏c��d�<��,��))_�)�U�3��7��sߢ�t�������eXL� �N�Iz���Ys�A�U�y��B�K� �"w��C�k���`r!��M��ϹXlxV61EB     400     180Q�1�B��0�y��$��q�V�O���l.$:'��uF&L(!�KZ
�ZM1��@����x/�o��I�i�E�SvD��)��q ��B��H
)L&�4vi��7����_���դ�X�[F��pxEΛ4�լ_0t�2��z`�qܧ#�������)�y�;��E�e�^q��)Qi����-5�����������Z��^�v�u��Z���l4���z��[K;f��0Կ���sDy�ȟ6>%�u�~��˓�۔W^H�Ƥ~v��>'�Vb4x�>���FC�ʁ��m0~�~t!�����6�5��:e�
����R���`bq�_Tn^z]邭K��`��	�a�;�G�����ėC������o��XlxV61EB     400     1507���*���{!��q�x�K�w<���jѻ�tx�N�$��Z_}�w��Yؑ+����Ӭ}>�	�y���;�Ck( ֌ ծצ��azжOxsU;�*)�e�H2X|���%�:��fU�sI���_��Q�*��|,�1t/MÑ^]�Ĩ���YVe�i����{l:�Y�5 �Q^�=��ҩ*/r������ǅ��)!
INw,�H���XVn��K+���i�*��(�6&����F���� ���t*�;�6XK��H�����a;8N�c��|A�ӛ�3⠹Cr�8#����n{����?s�|���j�]#O*�E���_(I�W�hVc����*XlxV61EB     400     180��������������\�-�6�m�@�䊥r�ޓ�`b��YKC���l��=����~�󶨎��ܧx� �o/�g��P����|�H�T?��-d�0T���e��b����uF8r��6����0	
<���65仁���s�L�~
U���[�]P`\�*��T-���4����\�?y7�6�}ƭ�"e�j>�l�pX���Z��W���j]�>}���P'd��J��G��pV�ъ�.�f$����BU;�B��궆��HjN㚗A��d�g�eB��isi����}�R�4K���;����s��)������$����������϶��6�@�R�o�����YR�ٙ�c��[۫>�s�W��vdk~XlxV61EB     400      f0g[�Mk�X�	l������E�gؽL����+��1�6����V������Z8]�Q +b��~�,�����,3�eM�	�s�7���H���W5)xF4�IK�Y�4�0>b�1m��N��!��:���	�t�j���וӝT-j���~��� G��}���=��N��s�&>��/��,K�bH�{��:�$_e����:���Z$�ʬ�L@�
�,%�iL��պF	�y1-�:�<{{��XlxV61EB     400     110�$z070/�h/O���.���O�3R�^�rUy+��L��a2�yϬ�
5��S8�c�֩��[/׫@*�,ث=K4�z��j)6�����E��t���8��og�z�����d{���h���s��#�دv���p��h5���V]�=�!N��{O�zIB����=<˥Ѿ��H?��s��� ���y˾�>�����@��/��d;��C�p�a���`�v��g��k��R�+{n�$6n���>'�����7�����{ҥf �vXlxV61EB     400      f0d�k{�ڰl>*X��OY.�6�0��p��X����\V��ɶ܏�49����)�d~�
��iMח��u��/��L��j�_<��C���P�M�7��*)�x�t�A�O�����o�j��w�%��� ���guzQ���Ҟ�Rb�9�zP���
5�;�%P���!�B	�>);}�X�Z���0�3���C�|�$>�aD��������#:D?1�������.ج��;%����e,�z�ZK�XlxV61EB     400      b0�2Ha_���{
�J�>RG:/����'�"�j=1��K, J�[�̰����=�H���z��ʧ�_�ߞ�s�&������L���~�<zَ�*GO =z���(��d�-�zW��x�i�G2	'd^�n�q k�iƓ�14�8�$�$�}�լ�Ѓ_�0U�"Z�1���ت�[GXlxV61EB     400      e0N}CXr�Hw�d?�4@;���l��,��R��K��A�J\U�5��)@���*�
b;\���1�ŐR~�S]�	%�-�Z*k/�89��������Y����3�v�	)��J�S*���.$�#d�ey���Y���cx�f4��or%�#<�~�	���N�k��<��$�c&@�$���}+��kh���ꏰ��N QX����EjL���K#�&?=��/A����oXlxV61EB     400     160ޯ>?�C��PF���x��J����)�1x��k��	B��x��G�&���>���ίm�kė;6�F���i2~2Br�>{}W�EG���S��OM�=BT0|��Xy�Ee�N�Ô�ƴݬ�!��+�|�k�Q���sk	1����3%�gq@7�����vRۡO"�1�PJ���#8[����<�#�7Az��[�^g��b��3�ǿ7��-�_�3��M����(_=LK����	u���aGᆺ>Br$�4�f��r ��	:����ELm4��N���J����.xbU��s�㡹�z�bQ섷�4��{��w+m3N;P��%�5�6�1¨A:�XlxV61EB     400     150��9��j��~}���ic'�,�6�:�ꦙM��#A�2"�d��d{5�8MrZ�e�h���H}�m^�Y���{��#m>�ú\c Gߖ�1V�����HU\:��m��[��ό}��֭���O  6��=G,.t�i.P�*�k�XAgw�59_��_��`�7\/�DL�0k�'�7t�ǕGU���ܜ�����:��7��c��S���{��C]�*�p a��<�K������F\�G���9A��It�vA]�:W@4�(шa�ƃ�����IV�R�?6.L(K�L$7G$�Ac9K��蓯�	���1·�;���Õ���vXlxV61EB     400     170����Q��3N�ޏ�4BuUGy�3{��k~��FX�w8����6k�iGk����K��%��{c ���nuk�=l��Z�baa��;9�tW��4�P�Q��X����A�.QK���<��֒�I�gN�ML��4�8��2V�1����Pcnl1hԢ4	بrpnv2B�l|g�FVT�h�l� j���=t4��q@�^����B:K�ٵXI��#i�\8U�D�.�@�v)�V?�Wg�1����Ӧ_���N���c���K��og�G �i��(��~Rya�^K��������{�MG�/�A=}Z8�cI��M��H�aDt���˕Q�U�t�u�U��xr#�9��mzﷳ�*AXlxV61EB     400     120Y\ȩ��<�ܣ��-DW���Ɋ?խLٝ�ώG��1�{+n(�W7�8��MƂ0u�.��/���� �8�I��jC���M���U���<�1 \�f�Ҵ�ξ,�ĜgN�Ub_�H
�%9�Ӕ1�MY��n#�V�u�%��p���:�9L$l}Q�)��-�̈́a�u��*T�
j���)�B5��X}6G�\��ý~�w��6'F�����G��%$Hr��S<ۉ,�F*a�u�����Ii#��@��s_=��o����EP��������XlxV61EB     400      e0!��`z,C��_}���M���凗5�.�񊣌����Yy6Qh{"��֝D�C�����@1�L����Om[s�Xᱎ��;/G>�� ���P��8��P%��G�"�C��/09�c>�&�j�(ƕ�v�@��\��>QkfTF�u*��ؑ�O�5��ψ�\�I=9<�Kݡ%\�-����\������,X�n����N�ݠݓ��;s�"}�~XlxV61EB     400     160����\o�TJ{�0�k'�?  ��_:go�j�Vů�u�u�ƕQ��,�̳*���@85�a�'��e%�m=��-����)��)�t�	�Qn��Zo?/X�؄1�ʒ�d�f��.Z(OМ(��լ T����L[�˦X'���tm�TpGt[����c"�nO�RL�'���^�&_Ӏ�~`}����[�� h� ���p��5����_����(8�H����ϬBԥ�Ǯ�$�fQ@�=U�7�D���1�[^b�
���~��q�|x�fu����-�G(� ^_0GًIe�ӏٝgEL<3�ci�R�wp����̋�����Ey�+�ӛڪ^�gʓ0�XlxV61EB     400     180�wj�=��
4<��R� ��K��dX�j��L�f��ֶqk/.�
��M>A��b���h���5��0-"� ��J�#�_��E��y�ا�:v�j�ol�{�}y{*�z�>���KC�&r;�Me,&~�yH�-K'��x�W���3�	�&�e��0�����nB\�J�Hp.:BF!ϊBmG��3�u�e�>ˮ���.�=;�i˩�O}s)F�y�N��x��FH��\n�:��\Z5S��ϫ�)��Wb}��x*|ؒ.�鍇�м$$���;���i�7-G?qҙe�IMJ[?��fZ�g����J2���\o�-��g���A1,'Ә�z�ѩK�0�ChԺM������B�#�ۯ0���	B|:��AZ#G�A�XlxV61EB     400     140;}/_�vK��h��/ʸ��}MD�f[\@gO!��V��O|��_�<�� ����h�
w�$�=���]2�`�r���T4�{ԁ��,c?���n��i/ݲ��>H�!��x\�{���_wŸ��L�ܼG#����_�1t���4��	������>��t��=[�y�&�;q!�mcP��O��Qh�*�Q=ʄ}h�?
���ٝ\Љ0�.����B(�x'���o�Uh (��s�fY�۫���<nq��t�B��p�ZQ��H�DͦD�Nܱ��(�N�"TN�|`xG*�5�mL0�oXXΓ	���`qs�~^gY�.��XlxV61EB     400     150�{��)F؛oT��:s:��  K�UUw�*�����(۰�KVM#��CXw[ՂY�mH�^�\y�;	O�Z��d�>Zm|�\���&����p�y�)��V�E��*d9U�Q�.[��3���h#z�bΈ�-)4�ҽGf���l�W�F=������,5�>����X
��@<�F�j��L�UW��r|

�3/i���5<���A��M��aa���w���H�J��y�j�d��̈���.<^�.�j�#kA�o���^G����í6���U�*��F)���*)�O�UN>���8<v}����Y�m��%8�K�?�w�꒳�^m�0XlxV61EB     400     140���3P9�(���G����CpӪ;�c�Tt�ߜ��-��$��'��1�q��?� �0	!y�-d�$+O�|v.�����#��,~��a_���#y��a�\��f ��C��+j��aoS�f⯴ɯ��G�L���������@��v�^9���悖CX����IDL
��}�Ҩ���0E��nL�D=�'8�%_�n'{��et#�Q�$����U�E֎�yT�i,�"���p�R��?�~�AAͷ���Y���嘱QRXv�ϒ�пr�kK����Bck��j�PY�z;ZtU����]���T�J��e9ۜ�}�*�XlxV61EB     400     140��h��&*�t;��!_�򗮀7D�v��!�[ĻH���GL�������윦1�|��"n�&�5P���N��S�8Q>E��=	�gc�����P��ݺ���D'1�y�|�hB���^��1�D?�M�'
ӽ��'�֤�E]�H�pL8�c�NK5�O`�:�[����&r'�ޡa�]�r3�>�Z�\�Ĳ��G�H��Gy��@�0�;�{����i�4�l>�7S��t��7���06�ܱ��~yZ��؆�ɇ*ڕ#�M�p��N�;�"@�C�]bC��(���Iڶ�$�.y�1J�O��e��\�X����6�y�a�"XlxV61EB     400     180�C���S����1��w�����rNȺX�Y��;bV.NV�E4{�G^!������
&'�_�\8��d��<	y����o��<ʹ�����cϚ|:lpa-7������p�%�L�S���w:j[_>��1Z������` ��[q���H��*��i�S��J�Z��`�2�g��N��+��(L�D��c��&i4P�u�w4Fr�Փ��rp!����A6������-n"`�;�QA���V,s��4~�rX)m�ĴѰq���QJ#�e� ��{�
̩�����X>;C����^�ݴ;�`�"�R�-.t�w��l�2%�`~��a���s*�9���d@�p��8��$��5.$O>� OIm�U�XlxV61EB     400     1b0W��E~yy�O���/�d01�u������~Ԍ�(%%�a_.��ϴ���?� ��q(F����{�W�fɵ��UxX�����2���� �Dy��_N�����#A ��_��"���H`}�I)�^�,��G�ur��d�e�L�� ��ҷ� �����$6v����($݅('�ҼS-�g�λi�ڈVi9T�D��Wp\-$�˫g%8�ʬ��]�9�dSCտ���ꎅX�v�F�j�cܧ��}�4��9?��*��� >��=�C�	5�R�Ө����*��^C��)��߁D��o�%:�u>����q�t<�) 6u ����d���v�L��9h��9RTSx�%]�?��'�2H��ݬ^��߸�G�:�s2�&�T�lY�Yl��F�" jG�����|51?�S^m�?�$�;Yx���XlxV61EB     400     1b0�V�CN�~Fi�=c(n/(	���휖�%�%4�ҽ֚,�^/N}��������� �p�����a�u��&�,z�k���D��Xa��VX%�[pk�;�����ܮ8�d���r�
������ƴ&��#�]�Hw40�5ߵ�X�C��M<014D.�,�7�=l�������'���	ꡬf+��LK�f٫�<�T���NۤXt�O�^���F�G}:�og�o�Т1L����V"\�\mjܚ�]+�$va�X�M����^�k���A,8ѐ��C5�	hl�\ta`����@��c���.��YW�t�T3�H1D�_���V�1��/��-֘@�@���ߠK86��*�/�0���H��C�q'�����f�脵]Y}�]����WI�/�t���g��X��"�I� ��t%�XlxV61EB     400     130��{����b�xO��C����J䵊��=(�le�&�=u��l�u�����h���#j`��ܴ �l�*ɭ�]�~���m�9MS8�aX[-Ճ�yr+���z��.�2�Z�Z��m�G�9���9qCj=n׸d��� �h�꿿]!��ƚ��E{~b�R����a=F jr��w?��<x*��g��J����g��	�(P��L��q���ޗ�t�,��.�x�W�[����K!<�[<F�L��e����������L��8�k�M��PQu��0�f(�Hƻ�
�F3E��XlxV61EB     400     130?�1	#�u��ܐ����3����u�u8�O�ǈq����TK��p}T"�>e�
?*�b�� ?,РR�<�/��r+��m���Lb�hg�s��Pכ생D4�СoF�S��NR��X����G l)W����*.�!�Y�\.2$��Q��\����#4s�N^-�U463��1�O�K����x���g���
Ih"Q���`�l��d�h��.����(�Z���y�	�tX�I�4�EѤ�p�����8P��($VKN�R�%����٨�L�e���?�OS��F��r���XlxV61EB     400     1d0�5�V��H&z^��ޛL=���~\��c�ĤZ�^���x�V�h�3o�ռ?'_�6����C̀�F�����`M!�?O3AC�.�"W��{(ŚF]F�0�+;'�c�[@������=���0���ļ�n�-OU���{�jV#������v<����˦�`E��Y�G��?����p�`�%.u�p[J���=�Bw�*v�v�L�3u��D/�9~��N�G�ǑEZ�\���N��o>��%mu�U�n���9����*.%�N�z�퓥<"����mߨN�S�njj�_uw����ː�q����CJ�� NrC[��T�;b$�*�|OD�g	�q'
k���M�v������G8A�1�6�0QYvqV�%:?Y�^ ��Hn�-*�K y9�	4��'�dŚ�GT7���]N�	1I����Z?E�yX�@)g���U)��XlxV61EB     400     110	� O-k����Yc�UO{0V������^���}7���'�G���Y�m�kf�~n5
�KX�\�a�!�R
Bj�D�%�bj[�̢��%��g����_��;M�V�ۛ`� �4d���k���(��Y?��Q[���$x1KN�������ҢI����ml�4'렆�����cow�z��q%�YINX���o
2'�ɗ�[x��շ��|�^�1� '�1�bM�����0-����u����n|"�u�	�E������h��XlxV61EB     400     110�M�+�q�B�%:n(��q`{����Q�s��V<��u�~��U�ㆉ���w��)^��a��?�k�g�g ���9*���5��O��^�<�j�m|�$?�)��/��j��V&_H|�{��H���&~� Љ��
�fa��*��sF��T����E �c��;j.��9�-M��nAgH�Cݫ8)�جN�Î�aҗ����u~l���X픈��O\��觃"��������1u��=)d[�� ^�,��Dh�[����$D�XlxV61EB     400      d0��pl�|����gTٯd�&Z��8c���;�e%z�lϯ1����o���F!��=O�*��0�^��o�#4����"����C�#���-)F(���a��e
�6�7��>j��n��k���[j�%����y̓�ɗ����,��F�s{g���,����S�f�����0oũ��K�J._է6�&��+���?��XlxV61EB     400     1a0�{��v�	��b��#<Y������ߜ��E9ʅ������g�����~����n9��*�UXBS�������%�\�a�
�'�2Tw���Յx.2�nX���Q��uwZ/8�;���jW���gGE�l�'M4,���2͔8����JH��G��޴���e�+��9$��b2iT`+�� ڃ�,&�P��@��_ץ�x"c�<��(!zwd��	8(��V9"��G�NX:0{���@�U���RF	�^�:�v�&�,nR9��d�����p�!6���7�9F���l�ڂ$<����M����l���3YE�_�}t#UD�zQdA;�=��Y~W��]~4��di�/����"U�V�@�����||�
��b���֯�������-P�bk�%;�
�^3����XlxV61EB     400     100\x��'�)r!��ˎ��0��^"�Z�K>�S����M�%y�߆�}7�k��=3��z�%T�gsu.=���L:\?ς��?K�L�N�����a��E��i(�A\�~��~D�τYK��_
�\�$~ʃ�$80���wт+�	�������<�doxƼ��eҺ��G��wJ���Z�UO�Q�� �>�JM[�G���1�G�M!�g��B��J��١I"��+ ��
.]�+U0��!�o��,=XlxV61EB     400     160:-��6����I;.�YrN��,S�#?@VT�����)�+�Tв�K j���^#��u�kRe�We��U"ޙ���FU�.��|兹�����ɑ4�E��b�;ޙ��$��3�#�>�͈�}$k ��~߹���m��YEkf.����У8o�g"�����.��j��R�+��Q\L�3P�Ij�h�k���ΧnL�8�k,���w,�������7d(���`��.��|�v* r��/z��o�| ��UV,/l+��SO�9��9I����a8�t'���3����i��;s�֥u�Am�	�w�y�����K�Ao�y�x�J+�ءs,xP*�D��[XlxV61EB     400     120?��[u�oٶHZ�*H/�u���k��zT���l�_��RZw��!r�1�$D��L2�}Η�GG'�! �Gt�4 ��,0��;y�I�l�0���i�Q�-��ntE2�P-��4@{q���V���	(Uv\��t%�FRܼ�b1}�UN�7$_٤Q}!����bK��W�T7��@�����E�+%�v�xS1���9v�!��j��7Z��&���Ar��U�9�|2��d��4QyF[��?{BP�`���Q���I�&� ��)G1�r���2�UXlxV61EB     400     1c0�o��S�^�	`$���8��W���
�8��^�P�](��T�	Ǟ�B-�B�(ΰ�b�X�K?������0��HB�it�ҡ��9ܪ���c� ���`h���olt�
J�%�ʮP��jo��]�{���CO`�ܖA�}�Ww
_3o6l!J/`9&;��m��B&��Ӌ>�^�*�vi����]�<yO�vN������=���Fn)�<�9��"y׌��_Cp2<#�<�'|��@�QJ��cCg1O�_�nV�K�����<A�D�7��h��L�S!u�9ֆ���p_k��p�'����[��s�ˎ�s�����R�
ךsQ\gt��d��
LB�(-q�:��}����8� z�N��X)��V��O��W����ҽ
28'��-�� 0���4�A��Z4�u�n
��@�9��Bؒ1}�t,!q���XlxV61EB      86      70s�K��]�� ��=��6$Ǌz��;�i�=~5?���^�����Ы�G�:�i��;	
���W�v'	� �³n�ד�K��R_���ɋ�y��~��f���n:�z�~