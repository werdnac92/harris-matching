XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190�Qs���I��B�{�c9W�
�^vJ������K�D sJ� ��4 O�L�7M��K3��a����_�B-i�@/@j���V����HD��2�����=`�b���e6	xu
�'Tho^��_V�0��%�'���3H3��/P/_D��"���6�(�8�V0����qƱ����V�<h_�eН���8�ѣFV��i��foW`a�v�_�sӯ�aܲ����������]��I6)_J��)T֯!�4D5O��g�G�hL���D$:�-�E?�ݠ��q���SP��� ���A�uD��زҏ� 8(!���l�	��<���nQ�p���!$��/��F�����1��;*n�>Xqf���x��Y�L��E�V���]���-���O6c�%^��/�(W����*�XlxV61EB     400     130�]C��0EWÄ�.+%I���s�yt�6�+B_����r�،z��N��A��4n�?\��m^wc�r����@��@�nY�57���v�1)���
UiD�jJ�ؓ<65U�_���l^˼��������=\�;{w���.5�;c)v�M�&	pq��Χ(H�ܵP�nD=�h���.�]&
@�CL��l6�����ܰYٻY�qx��&~c���%Q;#�S^Qw��ul�z|����9"���իsJjo���qX�:����7_��L�
���3Ȕ���fF9�룁XlxV61EB     400     110�F�
�%���B!(�</z��H��\��^�ZF�1=!8�Wܺ�Q�rO�_x����4���n�X�vֱ$��1d!�O�}�&�0x����f��!����������F`����ng��gׯ�������鎆��n� }|c�k�
N)�B���ᮟ�d�e��6����_��pZU#���:��Akj4]	0�I�F�d ���c�H�.Щ�T�*��	���Vۄ��C(�H7̃�$���1�w��0&��"J��p%�sQ�XlxV61EB     400      f0I�GG&����y_�	ܧ#^Q�K�Y��	����`��4:m����W��yu�eq=y�>�=�o�0��ד���C~�1�p5)^U�X�+�+�C,X�4K�R�Cs8�s�:�z���ξ�Y�b�,f�7
>F��@R�H��G����h/���"���[��F���z��s��z�//:����{��3���R��5�GJ��n/3(�fw
�R:-�h1m���ʌ��\^��U���̃nXlxV61EB     400      d0��SR�����i���q��]ݨw;��	�?E�M��Z�I�k�dz�pjFR�4�)����m,�xq�	%�� �7�m
,ۭɢA�9���O!~*�~���ـ+�d�j�����4$*����^�����.�=�ׂ�
��O+�����]���dѩ+'kӵE{��h�Sᴫ��[�ɫ�	&��`��c��*�o�R�XlxV61EB     400      e0_m�D���\V�9���~-�~����l<I�A/��l�[wf�(�τ�n@`�񷟫բے�Ա5{W�y��}^���B���.�)c��pg����@�4r�6�6P�P0��"l_H ;H�D#�K&d�R�];^�̖1�_�y�p�?������/Y���L�&�W������i^���X�FwD���&l	��.�Z�^���&A��kS=����&�[ߦO�k��0XlxV61EB     400      f0B���U��-}O~��FSü)�*9r)u��7�ɢі
����Z�r�q�*��Ͼ�<�� ��gZ����4t�&���*1��B�Ӣ��=�1�ǖo�A�"�n� )���0��
��:ӂ<J �+�gС���c�1��E��[�&�_��z>c��;�Q�j�8����YepE-���
;�
��4�?��W�>��4r�6b�p����Uds��r�?��i1��>��4r_K�i��XlxV61EB     400     190�k�:z��/������VX�p��<���n��8�����iǄ8��D�vG�R�w�hc��-D=4�<�;�A�)���'��#����L�ԿCC����)=
�6�������>8��Sqt�ژ�n��gtgY�+I�73����I�wp���f �#A�ȖV3�i|�[����Z4�db��?��L�=����Y�7c�~%�4�I�>��q��rH�ꉙֳDa)��24�_&�������A��Ju�Dn��"X���X�{ov�'K�,Fj�JVQK�͈�.���d@�9������_�	;G1�u�q		m L�2��`N�y/�)�6(N|rYap���F�h9\tpl��IQzcG�{�Z��-����͐{�c3��UJDXlxV61EB     400     160ʜ����Hg+����e=T,���=ZzY�##AX���ȅ;�:���%�;�7�$צ�#�#�{=�S�����5~����o%�e�M�`�sEk`�R�Xd㨟�Fڇ�?�m�P����X���T��^�Z��ݼ��~��T�l�.�x��k)�'v�ݮ��s�U?凱��3��ٵ [�5�gu�a�P;?�`o��A
i��%�d�����z��~܎�7c;"�:Z�6[Xz�d�ccPo�[~��W��F��`�D�(ӝE�a�c�IF"�
�2��10NfbO��X۵�V��<�!���߼���\Ѭ+\�m1dXj��gR"�����88Q�\k#҃x��XlxV61EB     400     110��P��t���V�L�2�~��W�����ۢo�	K��r�nu���C��q���l�b�^�?&�pR�jT���1���K{��K4�۫?q��G-V�Ä��h�%菊I�N�lE�;h%��#k���Cn�]�� �{4�d�/�"�;�LN����d��h(Y�d"G0��5"ҫǷ��v�%�㝚��U�p�r� 9�.�4*��+<̜-0B�@3#"�<s����L��f�M|?m����%�0����VʲT�bt����T�ifV�OXlxV61EB     400     150ɐ�/�:���ٳ��ą��aH��M�K���T
!@����ɟ�zH�on�S�8M�#�>U�V�\"�����.-[�^|
�WA�P�����u�^^�����H�9���5�CS�Vg{�؋��s���#�]����P�fb)~�{X�@&�b���!!$l�F���FKbj�g_�wK�Z5K5/Gp{=���{�N�p��#��Q�L���&�X���Mm;�z��_�j�4�$u��B���B�/&�i��YK��la�P?�s���`yW�YU�J�c��K�d1tB��,R�-�3{�H�j��kFs:	��������\u�o�7XlxV61EB     400     140�󖫗Vf-��f��W�(�����+�� +��B�tUV2-*�w`^")�c0U1's7g
m�H-�}�����n�`���X�&��y�O����FT�v�Y���w�:�R�@g��y^l��cX���,���1��7n!5�ޫ�'AБDH�H?��\b8�62m� 5�:[���'�rp$l:G)��3N��V^�>Mµ|T������j�����V���lx������y������H�Lr&p߱�C���g�w&��!Q��9T�4�f�<E����Zj�C)�!��Xm��d�ڏ�XlxV61EB     400     130f�Λ��\]	&ԓxy�S]]i�5���m�>��щ�&h��J	�f`�!�_7 !;�oEޱ&S�<��� ��v�o_u�(����{��A�،:�ۆ+�
!+/a�X"P��y�n����SאDb�{r����l��i���혅�쁡�l����!��L"{��a{u��F��C~�_3�Y���0�{�+Z����+Zŭ�����<�s�^Vx��s���3����'�bV�)R1�qlE�'�?4�<"�6���r�2��35��_�$���f`�e!�T`8�0[��![n�WtM����@o2j�Y���I�XlxV61EB     400     100�gt�3a!b�>�b*K��1^S�F7�Gy,��
�;9e���"��C�0S*��D&I�!�Y��>l|SMᴛ�Z ��ƥZ"?%�.��bS�Ւ����)���%�$,����j���ǆ������B�ZO���)�9�w�&�9�������s\~Vm��p���hɭjxuP����	�%��7qg����W�S�٩Ng�u]�Q�jێc~,�Qx�V%�y���j���HD���������6|\��XlxV61EB     400      e0Yl���~�-��
�����q�Ѱ�(ily�lD�����u*51�$���WB�#$B5>�:�fz�d�d����I��/O��쇾���������y�� +�h[b"b2����ؙt����3j
��
L�<Tو7����N;D���kԶ-�&ZEH8��A� ��W�}�]I�O�����+�(�f^��g-CIaSE��<�B�.����}w]�b-X�U�s�XlxV61EB     400     160�R��,���� ��1p�,�q�F�䇩V&�(f]�� 덗/'A���蠍K��.t296<.z�(b������,�)?���<�L/�ӏ���1x)����_@�Gm�SY�*dT0x��\��W|9?�A!M�0��dP"y��r�m,��^�yi�VW$b/�L_��6��R�\B	�Y9�Gw�k�����Ó$��32�0p�*�P��HD�IqX� �2�6� <�#3bm�8BRBE�򖬤���_��g�(6CƘ	^V���8mpHn�^�5�Rx���(~�+�B�1�5�JT�~�ԺEC�˾������|� �����E�o6�]�n�C���E�>�y 1y�̛����t�@X�W/vXlxV61EB     400      d0�����*�9 ����"����ĝY�����)�04���T �6� �!9U��sM�R6�8}R�������n�rN6D�Q��5��׋��_O`K��k'��,��k�U�g�lg�ϳ���oU�OS�U��X�҈�Y���р�W�ty��F�Br�88���վ�x��h��${�T�����)�2�v�$�l�j_XlxV61EB     400     120� U�m3щ�uu^ 8nr���>2�$�@�ƄCMZ��X̨�[#��#cA�{7j�^�@���,ٓs��ؚd;�D�re��$�E���IY3Ҷ_38�L�����΃��b�F��{�'T�\��vO36O,2g�n=���Ѝ�7�v7oY��4�k2�]� �h>�L�[�|��B ���i|<���:EfE�ѷ�XD�R��O�)Y�� ���刖��oHz5Nލ#g�ɪu�8��t�[Xi�.�[�����W7�$�)6N8%z7o�D�L\˃o��s���p�JkXlxV61EB     400      a0m6�<wi`�)���W�j�>�(8g��U�Q���O�&tD�]��p�$�����D�X�,����F�cN���o���|�l�'<z���"�*��C(���o�7ܜH�=њ���W�"�1��@<w�i��
J���(G�����������XlxV61EB     400     100U�0�$f��T��8]d�%�6d!"(�fx굙�7�w8Q<��J�{M"i����k��AH3\0��(�f그�w���8�{�����{,���d�Mzoa$�5$l�ADn��K����x,��$�^4�� ���2|~��e��P�_�@����jQ�DjW�M;�s��S��;��%�(,_��χ��N�"f�,� ��8�N��Q�+L�v� r�fG��CM��}�ae��V���3�
� �<^Q�S8�XlxV61EB     400      d0�i�$Ⱦ*������<�����-ut�$ڤ#���"�Ǹ��r�"���Y���t�t1Y�9TGй�#�|���삘Z��g�RF���ojy)�{%���|��+�tꖊH�mzS���VF܎���W6Tr�.}�������&q�+MP����F�ۯ�+�y���N-H[�W�u| эC�X�'C]饻SR�{mP(�~2ugDXlxV61EB     400     130B��iG���K�@s�-�{��֐���u�g�͂�r&��_������l`�'m��'�h֏L�]M��d�{iFm��%Z�%���{F��<F�g�h��˵n��P�[�ʉE�$�̓cVҕ��y�N�����_�� ���"��5�N����栔[I�B�,�j�;��*M6��o�m+n�iG�K�A�.��-\�g��n*X{S���cX��`\�`V�^����AX�N�{0��C[�?�]������t�-�ꭑ�M���s:
[�>Z���f9��	�`�,T����/ǈ�t5XlxV61EB     400     1b0���5\D-�Nh�%�sQ&)5���#�g��%�{���
���d9*������4	���ӛ�~{F3;�~��cKT5��Аp��7�p���z�j���9�Z_����⛮����2E�0�e\Π��Ր&�_b�B7�<��q���,mq�U�ʰ�|C6m�#��,�}�H��Q��A��Z�,*qqN�������⣀D,]�џ����EO��k�e�v`ʹοpi<���[݄�3@���j��ӿ�<�CÑDkc��2@�̠B��g��uk|f�V� 0gU	�ɴC��PjIleG&;�j'ݨ�jն~�	�f��&���h)G���tE 02c�i��CsUc������L�D[����K/��0ױeq��7��=L: +�Lo%Ņ�̳�&>=%�{������p}6%5 Wۏ�XlxV61EB     400     160lɎ�^9&C-�H1�A�.W_�ׂ�F�G�l^ZJ��F�w},5�c?�2MB^�?d�p��5�Ӝ	^<�!���ٴ��,ԉ�׵��9���RN[U�v�Vw�<0@GV���NJL"���JvRŪ��H��/�Θ��;'~� u�{�9!7X��tq��������w�H�����w>�A0�#26S��G��y~+zT/%��Z��O2�Se
�b���-Q˯�6r�gPJu��]�k�v��f{�Z�y�u����D�\r�X�I�r)�'�&��4Q�JT<��IFV:���6���r;�����`R{L�|����q�$��\F�w���{��]�AN�:mx��(��6x�XlxV61EB     400     1b0�q���"�����*�׸�#Ҹ�2�������[O�.2��1B�����~�yv0f��#�A��1f'�"���Ud4@���$�g'CE�n$*��<�3U������?��ܱO�	Xލ��L-
�z��==&�L�+ ��������Z�[��6��a�����9b�����EE8�3)��z:����Wd���
��%^�܁��|�+���W�U�|1�����˱�b;:�����"�.�=�7ŤSrJ�b�Fn���NO{�	��3Ϋ[	���O��j� 7ܘ�9w��S�KFg�y��:]*0K"�B��D������.v��µ�:Eyv�fD�h�S�{���U��X��`��:mE���N�{�#	�3�+81}u	l��H�gD�q�����_�����{Ư���\� ��3�w�XlxV61EB     400     1a0�8�?�m�t>"�o~�Pk�٧Pġ>��w����XN)�ζ�>9a��D _`��Rޓ���p����Țb=9_��l�\s�j7�>��ɇ����uz��i��kE���Y����s
�>v�X��Q̖��O)���U�dD�ԯ,s���s/H�q�����	k��t���i��g� ���-��hwz)�������۾;ڞd^W����4#=�\Z.��C���q�L�Gv�P0��I�i�So��2���L�
�~�6?�zUz�����%� ��p�E?���3
�3�����@��̰��̙p�U����:�aog�#����3`�-O	��}錐	�@mhb��S�Q���?jǹ'؋�;�I	Y1�� `���s����e�p�X�1g�،XlxV61EB     400     1a0t�L?����$�>#]��A��*
!Sã�ɭv� q�;�s��bb^�"���.n�4&1�$F"	�j+�!x?#B�%2Gޭ[Ŧ�OPYn	l�^@,�R����gT)7��6,	�|�A���Dޑ[ⲭ��{��������R���5X7�3�/H��P�y�u�\�sDFW�
h�ӫ�t��h�yfW� K ԚG@�G�)P�߀P���{�ݲ��0̘���Yi�Z8'�>Z��du�f^[$bL��G���p�N`���G�G4w�#�0�qS�]�U�R��m��t|5˃��yO@���:�HD�nQ���6Y ���K	g�x�I\ ��*���6o�?�<�^�"��(��ZG�[�� �)\���z(�t5��v�Qp7�k)d��!Uut�_���tXlxV61EB     400     170�� .�Oc*���IT������I�k����Z�ǷV����w�qto-C���w�s�?a�e��`�A�����E��tO-|��BK�fNw+;�W�d�67la ~{b]���n��쇉��7�BQ�Um	P6k�����I�v�Z�q���9h�6Tވ��_����q���l��S�2Qi�%O���K��A���dCu�5��F����Rύ�b=O�����!J0[�'G�l9��+�ֳJ3ÿ�qN㐰:ľ@�r]@����ǪO��m���K����?��~����>G���B�`b��;e[Au,{a������:EI��;���.h�|����4�ioL��T{���֨gi:�z�96�G��BqXlxV61EB     400     170X2��A�fC[�_�]��O/�C�Jb"�-R��ڲ���HDZZ����	��~����\�s�5t��n�]J�]��\�?�;oI�D3�pP�!JT;��H���=*@�g*�e�-��}���O
�q�-�a}��l�*Nfyr��:@��E�qU�t׼|�,@j�ϐ��`����)c�d-�B���Q����[{S�)�F.��x�&�*��P�=��,lbd���\�]��Hx��}�=��K�:>s�-�xWN074�%�"�*v`]�E~��߸�r�����m��d}��i��
*r%-H�\?��"P,[95��n?�.LM��=_li�5����&�
� ���M�����^�\lkn�����f�'XlxV61EB     400     100^I,Ww9B����_b��	2�~Ӛ�1=!���:9	�yD���.dXMV��5��I�z��лaYk29mM�W$��/ufZ�77����d��y�m����.0F�Ħj�>~���e��2.g����֣�a�x"��HL�.�Σ�AX�!����!�VƘ���r��(�M8����;���ٲe%�ЦV;�uiD���WEZ�eC��AJ�m�9L7����G��?<0��s"bx�n�Ps�O�
��XlxV61EB     400     1b0M�Y���i�N�8&8D�PjZ|�T����Y��#�X�/�慉�NR)�&jժG	�G� �4��߱S����;��|��D�O�f��_�9h2ae}fA>�6�}�އ	[��L*L�����!i0v�ԛ�|�
ۿ$��5����fK$F��!��w�8����kn��XˀNޒ�)l��*%���hb�1��� �m(����=i��n�i�B%#�Y&���<�>.��w�?͜��ʲA1`�D9���/lO-��T�i=z�w�Q�7]|�¾zև�wg����5�)hn�L�dPtB���!WNv��hTb-]�
6�lA��n�f����mm���OL�0�t{-��ǳ�q�]�E�������w����O�mJ����n���YU�<�WBZ�(XA�/��Ah�K���8�Ot��jrV�8��,�XlxV61EB     400     170~���y��k >�'sS�3"fI��&$a8�C�$� �*n�2ē���ٟ��i_Ӝ��.J��
-�h#E��EȈq;i ��r�t�a�N5��[~e��Q��
�y��R:�>��
鵽��>��٢{�y�:���;�z��R�y:Sn�*YK7�*x5#I�q������J7��5��NoN�U�.��{ȎsT.�څ�6��e���R_�5Vv��<,���1x��s�q�%���)�m7$>-�,��[�7�mx_�������e����'�{\H�A�������rl$�� k�		8Ħ�` �!F�f�!=�1+�S�%��i�2��vs4p���}�/�w�MY���� ��)|QXlxV61EB     400     1b0�聚��!���t��fWшܶ�R�[f,~ڈ�[e��G�fJ�o~+X�`�ą)+d<�u�������p�����x��ύ�/{?�-R�W�Q/2���$�L��;���Ah�~��.{��V��$�G��,c�4y�MoMV>�#7#�:|c_0�L�g�V�:���ϖ�]a��.(c�@�T}�nV�s�5be��VKYv�̽�[���Dn�g�.����,�HG�kM���-𺈁���OfY���y��t��7��CAZ��*I �����1W	��Q���~lѿ�E�1�]�`��cNN;j�t˳�0��r�5U>g���6��I��0c�<&[ʲ�rͯ�s���Ģ�VEf �����W������H��y�9Vi
���B]�.?�M�	x�m�����r@�_�nC�*L��U�X�XlxV61EB     400     1a0A(���6�ޑ(���N��9y�ǃ�P��j=���wF�2��YZ�r��f�@�x�Z���;��J `1?����*ܱ|A���y[RT�($P�6��B!�O�]E�}���aU�nE�_��R]	��"^�b���sIt>׹*K:���3�]�
~�����~� <�1�qxYə=��4C�ݯ�ۃ������3C2��ڗ���
/�u�5�x�\�n�67��|�Z��wE�K�WS�q$+� �i,A�Ub]�r]A��G��5x��2o�|�S�X��Ӧ"OKb.9<͐Li�?<�˦�Hv�YQ~����7���C�3�q��a��`��T��*l+c⡌,�e�נ���g_��P��2�p����JG�F����U��;�T�<���i����)wX�XlxV61EB     400     150��`V�$���~��Ɉ��G�<�B޾o��-��)�Bf]浥�ܾ��Q)`a�|u:`�a3|+���0�jn�Vo�6�4�0'����/!f�(%�6��uV��|H,})m^���'d�Gpɷٻ_��������P���K����@<ژ	��Ȥ����䀱��O�<�\�}B�ص�F�aod� xd����o)�YQS[h�֜5?�T$�����D,����.'o��>[��-��OZew�!q�N3/zs����Q4B��FB���S ��5��P��9K�1?��{j_劐��ݘ�{�h�>V�w���r���l��m{O���O��&ڋ�0;�XlxV61EB     400     190�BW�S���P}٩�����b�A8V��j�󕅔bO�,lZ�y{�����N���%�[r�)�*{?;����PT�yo�2[���*u?��q9��*v�oq�oi�in��uo����N\��n�ap�ZL���S�M��	�d�D�}���^�'J82D&�sA}"�Yǩ}�f�_K� ���ʹ4�9!�ݡ�	�>��%(6HD�J��zt_ ���[X�c��R�R>���ȲnB�}����E��L�_|̧���4{j�Q��:I�U-{��B�`Ow_�!���L��]����D�e�'��bj�"|u����MS��yo�qlB�~QA#M]󏬼�É�����7������jT)IR��G������ajM��X]Z"���a��d���]XlxV61EB     400     1905愈EL۸Cȗ����TC�3�b3��{� �^�]C�0 L\Z�������:��i���,N��$Y�\���V����?CX�։�n�O-@DM,�Xer��;�����L��m�N� c,�&��E�Yo4�L�%z]�.���:��`�_`�H9���䓪6��_)KA#M=���i� a8!��I7�^K�a��w��c�a0�v+�[%%،!��P���/K�l��bb�����ď ��Ɇ�X5KE�7�E�:T�C��b/�TM��y���S��$�ĎdVn���$����!x#������O��޺M�m�v�4�:��;10�2�孇�ۜ���&�A��B'��y�����Ub�;zy�Gq.O�
O͎��6��`7���퓥c�.XlxV61EB     400     190��l��-��:��^��E�U���n�2hk!��M����Y���7Z���&�5Xm�B�53���5�Fƕ�gU9e=��?�j~�x��:N�a��3�p5xFk>OZ.�9�N�~Cu��(=\�%���(���9�j��0�]Joi���|΃i�$�q�YW����G�豈�-E{�U�XC��Ovad���`r7�N�4�~�%%�����4����3p}иap��Q�l�F�B=T��K��_�W����Jb�Hl*�Dމ~������Ʒ�U�`q5���KZ]
���#��i`V�܃�넫��J";f��H�o�2ir;9�K=h[����e��9��>)��E#0ͭ����I�0���� .^�0�>�¿:�'0=���UUXlxV61EB     400     100(�9�LVb���ʾ�5����3H��*�P�J<�M�.����d�l?�ȧ��u�� �/2���đ�L<��Q.���7��������ERo5N/�,����7���a/�cx��d+��3h/'/7����Az����+�^�j���1��[ڽ& [b��Z�9��A���4�	K#�|���5�.�^x�U��S|)��N&D��L|��l�`6;l���4R����8���|u�S8s�S��Xĩ�w���:�XlxV61EB     400     150�Cac���O8�f��]å��VGp�7Q&Sh��jo%z��]�J������1���W2)U�i��r�U���.G��7��
�lV(�'$����d�%�l�U�LO�������l�,5MrxX��M*;��E�#��߬.����-yۚ�&w�\Vj!��6��*r�tu���]Nή�a�v�����?v-��.	���Ugɗ��2@�H����$�����,�����{&-��L%GǮx%�nňR������0��,�LK\W�c���G!%� R����[���0(7=]���k���A֚���F�i!jm�@�`
��2�0��}XlxV61EB     400     120��D�^֬�sl�5k�|8�D�����&��331�f4�l��u�%c(ʗ�e���Y��뗿?�-p��p,���P𾰱�Vp(��0���sK9���wƝ햖���[Jͅ9�ۡ �0�������	���Y�=m� 	���h����I�}V��U���e�@]!ƖY���:�=8Q���ڄ���1�.{��L�6�Pѝ9����#SH&��U�y�ݯ�R��'J��T��BX�)���Q�$����j�xN�uO��0O��9*5#� #� *o�3�-ň_XlxV61EB     400     160.��9�QT,ZY3�H|���AS�+O���e]�ŕ�o;Y�_~,�* ���}{;��B�s�jk����ۡ:ܢ2r�t�+鹸\)v�MI�h��+8����~R!Sn��Rַ��O,�;���]���.�z�ٞ�*4m ���`��H)}깑��P�W�h��W\�8HT�Z����?������r�J*ɳ������+��^�[c��k��j��=b�V�����>���a#~'o��U����e��$�fqƈih�"u��G�5#���i�q�D���U$�Ƣ@m�lJ��݋Uˊ���84�9���[l�ߖXXo&�ߖ�?�>%�l��d�nn�w�XlxV61EB     400     140=�t������R�(*1@�T=0W.1I�9�ꦿv�e�.`m���}�E��ڸ�Ų������q�|�/R�q�|�)ӱ[��%�B��4}��K��Wn�YC<Ɏ �t�W��t������F�/�y��VYz?Op��p4-3�^}r-wB� &"x����ɛ�P�����n�<�;���%�ŝ����/[��=Ub��	4���ohݚ���¿�4�߶���~��Uuy`E ��"և֦^	 ��������^����rm�A���4���%��upT��ž�So�D��^���!"�*TO���h�e��y-^� "XlxV61EB     400     140��5��]��q!�Zfj����oH<�6uV&]T:^�y���B)�~��_1���8ƽ��ӎ������3�K��W7�	�p�_j�l�$�:�*��$�I�J�*�D��t��V���3�#L�"�ƶ�Z"����Q��@/;�J=4�֣*p��
i��80A?�����"��+FZ� �,�s�y9/��-&����5�e����27O�V_�[�?�~u��e[2 &�{a�8�R*<�gh3J&��`RU��u��LTȚ�s���-L����ٞ���ʭ�*��#a�Bl�R����oRXlxV61EB     400     170���Q[Zz,an�����?~���/����=�9�be�e����nu'a�U�V�_v�ͪ���GZI�'�6
noc��9E�|x[����Qp���r<ȈQު ,��u���#�kC)��zo��������'��m�n�I��pU�xP��yt��Z-�fk<�.�l�L�X�%��:���Rk�&�u���ŽSX6���@����&�3�f�HӰ]�j>N��a����Мƒ���������$$����B�W�g*�2ފ���`���2X|�}�O��Y�|�++x^%T��^��7d/�!�v�}ư(�IH&����)��8���:1�)�I�>�OR�J���K��,��d����h��F�fPXlxV61EB     400     1a0N�����I�0��8�):�b��2��;6� vsa�Hz9-+��rw,�p�����}�k?h�ˠ{�)��\�>o�`,��E%ϼ�iQ����&=V�YP�X����c?�<?O��0� ��m|�����W&7������U�JS�v����5NE�:�q��\�i;u�'��O�U?��Fu+|�ah�q*��֋i�D�Y��l��'}�s;��g���v�Su�7l���v�A����]FNB�kj�Gi��qh�k��u�4��/��6WKB�Uso�~|����a��� �*߮ ��M��A�k[x���!�EK<N?�\��P��0�����Q���Wz�:�ǌQ���ԁˁM�
w91�|Ѥ���m]���rYN�M�Lj�e�Z>���Έ���n�q-.��Fߵ�%��XlxV61EB     400     190k)���&t�'�$��/Ob��
U����Z�{�S�'a��F���g1�� O��4vex�o�	_"
[OS�Q$&�	fCS����� ϴ0ɛ�EX��Ɠ�6���t����൨�&΂Y���yZ�=)�M��xi���N2`�2z_�1� 	ӌ��b�{m���1u= w�>i���l3�I��3c�wxfd�K�.x����"!W�8:TG��-�3�GS�O��hU����r�� o=]&��9c��#3lz7u���w�߷��B@ _-l2O
����
�^(���K֮	��z��ʁ�T�xv�+��lc�3]����L�x�b	`�]������=���N��>�)���fv�%�s0��7H Ѻ��[��1&t�=��{4XlxV61EB     400     1c0�1-9�!-,�#���Srr��;���mS��z}ǋ��:�~F
�� �!��V��D��ឈ���z8`����h��՜�z��M"�`�#1}6���y���A�1 ���	4���Hx3,O��D�>)�?8�ϒ�j[���&.��]�$.B�ϵ��Kn�` ���K�*f������b�iH_g�i�qjS-@2m�����e��D���t�˫q�
$��;����̴=��PS@�c Э��T*��c�c
�#�0P�c�SV���H�6x����$�w��ۑ5�QM�>=-��b�WJǰ�\W��W����ӜF�f5-�nDjo���*c��d��~��� 	�C���P�9Kڄ�S��/`�ҩ�����pu��HKWL@R��jl�����������A��{+�h^3���'���M13Ѫ}��t��l� .`�yI)[XlxV61EB     380     1a0�\�YO��^��T�VgĒٽ^@�v����2�Dhs�!Q����'�Z��i��m�����qi٩�:�|�+��K�g.�2�a�4�=�f�ux�<�&=���I��ͦXh�A� �[��o\�����ĝ���,藥���Vy�G�5�"�^���[����$3�r"Z��i1[�š�2�x�^�>T`G�Q�Ē�Ϭ'��T�):��:�g�H��$�[:]'�l�d�R��L��:Ĥ���.�gū��-!F��<��m2���6��ƌ���`��|9"�r#d37~���`�'�MS����3�	����ww�@>`�)X���L��"	��c�p���Q�0�%P�2�u���%<��݇.�������n�I�BZg�|�%��U,5ԙ�r����\Uc�ny��^�