XlxV61EB     400     140�E�e�?UW�����5����F(-R��&m��ٲX��nZ5�Pr���?��'7p�k23���T)����I0q�@��Y�5,r�~ع�E���$��2�<�XPF����*���e����>���z�*q��&4,0�q'e�IWU8��F.����*���)�!047�͢�w*��6�f/l��&�$�!����L'���&�V�N�����2W�"Q�kFW�3}�Wz��a�<��׺&M|ߵ���·~��y�i
�	��O�]��������)������Ƭ�TL�uC�ҷ	�1������`�=E(��-<8tn�XlxV61EB     400     150u�4G���h �;��H�NY�0� e�q0�fV{���A>�� j~���*X*zЦT�I�=�%5����g�vv�p��4���?�"�w(��.���`�]�<o��U����{'\p_XK�i;[�h�F�;�;!�А��ԧ�ApjLWG�	R�j��n%�^�.�g/*�CgT�b�K�b���{:�!�̸�Qr
�o�bpف��K7>�`w�ن$��A˭-�G0JE���]K��፱�L�Ѥ8.jK��|d ,*R�o��g,��Ԇ�[�P'A��_�Č�<!.d�B�jhbx4��8����J)�;����C����a�4��զDXlxV61EB     400     150[���a�.��9����?�Dg�N?lnA2`�	�:Y7M{�!�(cELS!.Xri?W�������79�	�(���VNGh͒�~�5����oX��!�9� ؛��ˠ��
�u�l������,��	�g���U=I���q��?�$_�Jb?r��w��c��]�A�S�~���V��9�;�N�)� �駄�Nln�p������m7�&VWد.���Ka%�J&�&�:I6f�uxU���Yω��A����sV��xx`R5j\,*�;�x4�������K�`L�]��U��i���~}P6���Uh�U7�呭�7|�ܔ9k>�XlxV61EB     400     180.Ǔ[�kv=5&h7�����f���	χ%���������9<��ے�Ix��Rޏ�̹��7�E�W�(ke?QB>�r�L�����Q�Ѣ�b_�i�ag�kt��	��B�F��Edռ�3ۢHP�D��o�<xێiE�I�&p���I,�� �$���yz&��7��w����U��4��/���N�
 r/I����R4
����K'��CY�{����骧�D�g����NȒ��;�8�J���¦��a�У ��UV*>F���7ya��/L�ps�D��W�dī�C�Sxv-
`�P���E��R��g��Io��˄�u}�_�q��2{�YoyBk��+�jՄ��I�y�Lŉ���(:ly��}3[}�e�%#|(XlxV61EB     400     140�=ׁ��;�7�_�=�r�7sP������uk�h�pV�ɅJ��E@���1��Kg}=xl�YS�#���Cy$�D���o��́��`�(�uV���]8oի6�P�n��&�[�<"�_��U��TE�a�+����xv�I�n[���ũ�L�����<�2qs��T�aq'g�Z��s/��	w�N�LUm�����33�' @.ihX|��7=�l��JzZ�'�t�����Y��<[:Uu�	m�cv�u�G�3�kȍ[l�h�*����B[ۤ���h�ˮ��`�E�(������L�` ��L����xA��:}�/E��XlxV61EB     18e      c0C�x� �RHi !W����r5fD"��`I��td�'���,�>YyTVׇ|��?�yp;Q�?y�����@����$�^��ZV�o��Z���� G���0+2J/M�s�|��AP��YG� t/�L�í�܍"�����-�S0���j�7\8t�ݗxM$��d�BݘIH�Dx�l:ӮCoQ���,]d�