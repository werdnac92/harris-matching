XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     140���<&45�܆��>/�Y�.5*���pNlń�/
�%�j#]Z~]���)�tI~�y'e+�K��mͭ��$P��xN:v"�R��d>�-���GI�[a��p�F	tpD��|<��		�y��R+�N(��z���=;��#�7ʯ�G��-��S��Q�ξ7K��b��b(�Z
��
�/\D�t"��K2~�K�b�����ړ#�x4�V�0��$����)�)J(���:ɒ��kVPD�6o�J��
r
��"��T�HS��O=C`mӭ�xK)!%�䎋~�.��ʨ����@��G���&8o��|@XlxV61EB     400     1a0qOU()p8�e3���G���	�
���� f� �b:Z�s����6�Z��t�8;�
^GW�۫��Ho�r�U���I�U��IO8͠�2�E3`���1Q�H�w+�J|ê�|��=�f��3_q[��\�lL��=ǹ�W���	!��LƌF�n���� !%��J5�6��>^,>~ob
�kK`͠�~��V��q�'N�����iH�%V��8�e�⮍ZL��X~���U�+�S�^�(�,��JA`���χ�P�Wsg���-��nײ�JaiS����oC�&J3h{�
ZH���.�L@5�@�7ċ+�("=ةӯ�]���Z���6?:���d��S�����ZG ��L��
\w�� ��ܵ8��$e��]������T��a�y_;͸T`�ϼ"0ܿX�hXlxV61EB     400     180�����%�c��1���os7T(�r���5N\�V8�2oS���*q򾅣	2�w_�v&�Q<�V���jF�cž�S8��6�-�~�Bꠀ��DM���[�ǃ���@�J��Q�R�D�{[.%���^9Ѐ�/,� ����f��֤m�u �P�Z���"L����E�/ 5sU���w��;����r�s���qC��)-/T)���o$屭�/"$�Ƥ�p%�$�.�U�O��`J�g�ql^(���	h�>ϵP�oxǧ3����T�Meװ.	��x�ƽ.F�"^��l������������o@ ��W>�tu�N������1��k�����i��Y	. ;�3���L%�h��
�w����>H��/�7��XlxV61EB     400     120��>��<YV=�X�s�敤��ٻ��D���1X;}���X�H���o���M�)za�ְ����n�E�2�^'�J;�s�ُ�ˇW�7���>(
�|�"��=C�bP�/
ys�g��i�ɽ/��ԋRu��i�ez�?��<v�l�F��mⵡ(�n�/_��"�d~u��U��J|�ް�h�)kFIH�G�d�/$������&*
Ph��ί�]wk�ǝ�����~��R|�R�gH��ծ�<:�)Os�YxY+.�	06;�=��KC���|���tU��*W���XlxV61EB     400     110}�G�� TPQn�b�E���2؝uoE�"i�!�!��枳rVY��
��b�]Z$�����rɼ��8ރ{K��Cdǭ	�9�+�bJ�� ������/Xa�F��i����þ`#��kf����E�i>��.��m�D2�C����A9��&�I7+�[ru�d�Yf݋�����q8�^uA�~P"ùU��d�*���f澮��`NX�8�b�����mùH�r[�IQ|�:��p��3��f��[@��YG�*z�)�cԞ�qXlxV61EB     157      a0�����V�=a�h[��;K�0X�Ͽ�4��k����T���l������5zι��4���R�h�1.�y����l;0��>���?�|���!����]�خ:����,z��[��HY��~�6��jbT)���V
nz\��E����uG�����,m��fb