XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     1a0�7�?�&��9��q�f4R�
8�����}�l���X��GW��A��ib�9`�	v�?��[[+wo�A��
���`F��,�g.���}��]���p�W�<�,>X�>4�y���������p'f-�Ν�Q���x6H�,Z}��а�%������h6<[}��۰C�u?�'�v�ƽ	�I���o��e*0'eF;}��|�2�ſ�L�^C+��n�qL��.}D ������a����1d���4o��.���B��c�E��j^��	��}�tĤ�u'�a�@�~k,�D���a���x�(F/��4yv%�Y0|���ύ���Wf�lz��3V1���nU-%(l�ӄT�rM�\��;��� 3}a~:Pz�R;�.�e �a�ʍ����3�fŮ�LXA*��}3f�?H����XlxV61EB     400     1808-Q�o��7��r[�S�N�E]j�ZQd�(n�;�K�&�zZ[�wkt��D/J�adt3��,��r��ˢ�bμ�*�$��@�7�$�����W���[L(B%�pt^��%�.:�t	0z
�ʴ[YLp����cQD�ቬ��blD��|�lR��+=�z�+��5c�E��у�:���о�l����u��|��ޣ�*O��`�)��ž�O�q�d�v�Br._�j�.��M̣^���N�e��;�@����a�;i@��p���[~�B�E*�=�wwl�H%H.�/AP�HXN7��5����-ʚNs]���d+�s�����Xu�߽�	R�pV	^���`���x��A���؏�@��o��wO���É"��q�XlxV61EB     400     170��ڄN��b�R��"�>ye��R�ЌDT�ȁ���撙Ts-���ߨ@5�T�8^|�aXY�	��l�+!af5�Ҫ��{��²Ĉ0sUů6(��e#��?��G�DU&cvz�켍,��pQ��#�u$
e�/����0N`��Mo�����B����� �{�K��h�I��%�!'%�XP�E$J,��á����m�$���+��O��3?4D�#e0�%���~j�mY�A�<J��RsF�h���( ��71�Woc'�;D��*(�3�*%6м<�D���0��n)�
����}"���Ȱ��7��g�K0 ���r���Ȅ�C�ϗ�z�n�u������y 8��!�XlxV61EB     400     1d0-J��B.����B 3��,��Z�$�{s�nс�2�}t�+�ys���w˲���#H�NLD�~%;?�[f晒�t�S_?i�,�)]]?��x�'s+=�W��?�	�P���8��^hq�G ��t��:e)~����]~��Z�Z�G�Af��wql�E�#,Tp
����h����U�ir�d��P
H�F}':��>�W1!�Jw�B�*��|3޽W$��0�g��) 4`py`,��!�Z����Vh��Z�٭`n�R��3��B��7���n��2��	���� �-;�4Y"�7h��o{+�j���L���U��'�r�8QV.���q���p���ۗ~?'U;]�����ԓ�X����lm�F�Ɖ�.zQ��w�3���������	S� ��%!�xj��*�,-t���j�WW-�*�꟦�����cj�Ǉ{�����(T;]�6#ԫT��p�E#\�XlxV61EB     400     140OsO<]�b.CM�zu�.��_�'�->(���qg�����H&���|�8s�\�!WC�BVɈS�1&�Qo�]���Y�W	�А�� g;
�x�h�;v�~f�p���6���6wݫ��'�����]:�Љ�4ȸ]�~�C쪖��LG��FPk����N�)O���
�PA_���Fc(^��m��h�2OA�x��V�ݷؔ0��m�d�%��xe$�58 ZƟUn�pd�K�YY��J#�������f�_�-ؓ�A�s'>��sh�*Y3p6�	�o�lh��z�O]*����tecg��2��XlxV61EB     400     1d0���îR�C�L魈V	x �&1�R?h�j��z@������w�9�J6G1��ɈG��Pߙ;u���d �����d��
gx$4[�$�"ָ9
y�0^����c�Ƃ�B��"�}k��N�*��^>�������b|5� �P.'6�Սj��j�L
� �g�U*��q�`T7e�k[�z��!z�3��|�?���ҩ1/��B#�I��� �'E��͉�V�#UP�헆&5\@�ǯ2'�bh�:яm�Zr��%��4�m�G�wY��a?K�.����<�⽃�sH�;[�.^~T�d*�<�S�"�ȥ.<�ɦ:9��O���
�pNki/މ�
�0KGU�3e'�~�x���ŝ�ʕH�=ǲ�o� D�]&m3xY:�[���!�+�.�������@�~�i��oM�cy�RK'�|�d�\u6R��2�c�uhTWZ��j3q(�.8�ny����L�t���G(�XlxV61EB     400     130�7e-��?B���b���2XZF��*z&x��aX��&��?����%��p�x��؊}l1� ��B�e/(��:w�&Ћы�U�{��G�QI#Ħ��~I�c����/�����D������E�xB�e�E�qٳt�&f����Z�.+�C��s�`�c�Ct
n-hN8T��a��D�I2�6���z�C���!ܑ�)�cz��#{ҸT"Q���f�Z+��љ�&�W�����C?d?6���6�U`�0��8��F9����_�U��q'Y{��I����7�,�,M�h��
x<6p}7�LL��vXlxV61EB     400     140���r�u�����ހ�[v�f�۟˲��H6�!x)�]��}�xzK����ladw�/�m�P$˜U�8�������Λ��P�q_�\��y��P���n밼�Tv�|P:���(p�"�#X�6xQ�>N�z.��nܒ4DO����k�OBR- �6bo	�ū���&��f�+��&O�:B�bhx'�Az���OU]d�<��M��Y���J}Რ�dZM���^��.Q�=�-�c;������@��|�#���1
�{�u�Q�'�i����|��	Ϊii59i#�g���T~b;��ڕ� @4�q*4���Wu�^5]O��XlxV61EB     400     1b0�|
m���k�����Be�:s���u�~A}iݓyJNn��pq%����3b@�!
���r���+;�+���T�Q�>��!����r��W˜��Q�q��<d|�'���gKY_�\����.1�c�E����+����u���#ꃉ��,i�e��;.�d����YW��U��B�1k������;�Əp'�0T�
U�ZB�pS�C�{��rb�c.}6QsH����.L�c��¹K��pc^����'b��IS�w�O���C��ݨHT���vSEӾ�8r�P�oO�+�2�g�hw5,��:���ݟ�t|�'�n�5�	,��N�실B��7���^���{��sU�]A6'�).z��ٙ�X]�M���y�'�-��U�k�"NB ���	^Q��Xf��<���D�C���XlxV61EB     400     140cr�1h0��zE��2ylB��2u�N�0�L�	��/��F�s ����V��%u��o�
m	��He������{���BK[�:�$��z���8KV$)�x4Ò�M�����u"�(������j8� �nt�x��V,'K��M�VqI�??*d�:�}L���:ǆNR�̻c� ���z�U�� M��Q��/ɿ`���"�� =z�okِ�����j�[��e��d�,<�PDeqt��t�]�b�-�T�|�MN�<�7^� �NC)u�OY��~z?�h:�Gss;�K��`_O��j��;������JJ��XlxV61EB     400     1a0���u��n��4�;�<�>h�Ӊ���x������
93�NȘ�pt�[���0�Ee�O ����K.���}x�1-���:$�8n�-� ˷%	���c[o������7���E�!@w'ŗ}WI[k�s���fSk��S�|�;�ؙUD���[Qx;�!��b����b�<ߝj��bC���C�f��s.��&�9.L���p�G-��e@˺�Gjʖ��6�ڽZ�H!&H��
|ڐ�nn0ܲ�R4��:��Ev������'f��}M�^��LV�w�X� �x���v����-�.�{Al/����My�Qh��#�B�ɶ�,]�
�h�/�%n%F�Wm���D�4nr_����Ж7Q����W�]�Ľ�؇�L�o.�3靤�'(�V�I�]�q`��2��.p��*İXlxV61EB     400     160_�[,�Ń�����W�vob|B;�Qg���d�/�P�5C�0���K���|P���QD�[��N�� �.i
'�1���)��(V�:�55� Du� Z?����[���ˈ/�˔�KoO�ټ��&����i�.����xB]9��h�������Q��
m�MxO��Јq!~���-�ۄL}�f9SJ�ǭS7�v����Qf�`%� �r-�y�tP"��Su�i�}���	wr[|2�?�Ro fh�';T��'DA�'8]�,D�nKu�Qi���U!��:.����k��Ej��8��A�J�'�l���*W�	wAY2�Bp�����$g{3�R��L�n�9[XlxV61EB     400     190]e�1�����+�+�������E4�Ꞥ�;�ѷ-���7[wخ\����щL�:�7���- �)	N��ݟ�H�|
�"�L���������W�t��ޛ��^�R�@w�~�2 +?�=���U�)�=�64�$���s�!bJ*�j,\�v�ɔ`����=0�}�C\i���t'Q��H����(�dB����[�^�q���[R&�ARMU��j��7^����Qo.e+��t�f�y"{�o���<�P��g!� ڢ�����,�Qٍ=x�iȮ���G�\ ����Rl�#H��D��	��M)L��0A�C5�.��.�&A����{�Y];�zi�]Y(r躐�q�;�k�j��w|��H�,���Q�<p�8l�1��_70R���XlxV61EB     400     190u�^DX�6���6u4M3�����wq����%:��Z�(Ih�4�4�\*J�j�.#.O�k��#n����%)
֮�9�f[�/0�]�k�ޘfB���&�� "L
����b@����W�\��ĥ`Y�C�#��~��;翄H/��_R��a���a~��D����G�S����s5
Q��p{K~`K�6Y��?����Z�w�8&�5�/d�Un��}����yN�R͇��B}jk� ~��lۢ��9�%�]��s-��Z��qfG�W�)*Oz��m1�Ƴqv�Β䌆EÐZqqB$�s�	5�E�-.� 2�ca�3��Q��:�����hfT[�Yjt����=�����p��F��~p��j�@އg9*�A���t�q?�RXlxV61EB     400     130���r�u�����ހ�[��#�	�qW����3����P;ɹ�!�v��Ŵ�4��4MQ�Ʊ�l�ɟ�RsԶ�,���#�2Pj:��j��L^>��5���F� ���J��4�/!k����OT�j���Bk��l�t��׶@7KL8���9;���u�1���g~V���x���`b,��VX7,#���	�mW�
�*w�L�]��_����gĝyF3M���T�7Y����cL�ո!f��-��Oj�d�b��X9�/�#J��;�[0��ǐ����]���'E�����!���]�}���XlxV61EB     400     180�Fs^�Z#���tF����$f�4��k;�ɩ��gHS�vj�(^�����L���b��Y�~[?��K?T(�)Ѷ%^����r�
]�%�n�� ��J�%1ұ&��Z�������y0*oq�T�M�f04g�w��O��W��dot�?F-<?�B͙@P�2l����z�@�ِ��9t�`�j�.��-��X� �[uIr��@J�����#6G���-���$����^%#�d���C�qp���K�.����5��M�q��Rm=�x�NwD��>I&��)_� m���ȿ
����|`��(�UhK�Y���$���T�BcCú,_�R �p��mv6����dN)��sFXY���q�LHғXlxV61EB     400     170i@g5�kK,ίq-{G,^� �r��#l�h �]Ȥ��q�B>#Z��Yi#��"��4��|Y��&XP�
(��Al�&�3�o�N����pf���n?��ԏk�Ox%�7T���4��PNd�[�z�mC-z��$�]bs~U{�H��Y��$��`�ɟ{�Y_�,��عb&��Ŀ�#i�!R����ѸX�N4L��,l��0�Dg����-:@�U4��Q�̌�fE�qD�A)������4�ucI���4g��S�i��/�2^�-���C� ��H�.��ٵ���n8���� ����k��`�۵���iE�c�;��-o����E�?zjr�!� o���kK��{89�a�_���ʡ XlxV61EB      6c      50(�W��Y�wZR�,�ޑ�2�2�<c�K�+2�}H�O�`L��� �)"���3š|1�g��5��Rmm�?8z���15