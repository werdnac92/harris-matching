XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     140�V���Ӏ5Ͼ�2u�= �u��:�e( <E(����������#Vt�jZ�'�G9�-��Mt�b�����٥������|�iǒ�}�W�S��8�t�O��?<=��6��u�j��[��@��D���ћ@���{,u��f�JFU�t'd�x����J:�zχ�O�%�w|�V0� �W�eM-Ǟ/�7^YID�n��}�6���q���t'U��.1>q�d��,��`���
�dJ��#=�.�YTQ6MB���l��^��R�,D���o�[����hg��6���NeV�Ј�$�mç�Z������A3����$:\�F�nXlxV61EB     400      f0
:Q����gR�U���`�E��X����pH��\�!5�Bzz�dz�a@�����'�C��H'Ź��!��W^�<�񼏩�g��W��9ٶO�.n@k������d���f�� )��,�aX�EB:�%���|F5E;Z�+~A��|+���?
�G��T��.�J�P�wVm�>��~��
z���2�R��>�Hf�{��.2��JLrn�
2�63L=
�
]Z���sч$� XlxV61EB     400     160���܂��ϣ��[����7�?V#E��St�'�׺55���-Z�כQ�i��&V�yn�׬��־]��Ū��q^[�
�e4��V�"�j��}d�r��q�|7���=q���X�#��:�w���"���qY�%'��(��u!��_�鐡n����]�*8��֓dl��1��gLK���`H�+�(��`�f��@��S��xP���R��9��t��k����]�̜�3��(��m�U��]�`<�@�ӿ��z,��o���O�@��$�<�ֻ�ćt~w�-��6�Z����Ml�t	���9t�}�s�&`�����ű���6�aZ�'��>�Xڔ3 B�XlxV61EB     400     120e����o�$ג����1#	oGpu=�@`=���ɟ�[��!��d����E���O�XO�ޟ�j6j���)�l�-��ꃚOT�5O@�]��`��v)�����R�ާ�
6�y�W�XQ��P�v ��F�+�CIP�l��v�:<��1ո��~f�����^�1�;���Ѱ9` ������g�0���^yz��^i%ܒ�#��P����;nIg����5Os8��>�T�Ǟ��G�X�����	?� p��K��ln����K+bl��u1b��´8n�}��XlxV61EB     287     110��!�u�I�}aE�2�e��d$*jM��n��SB��)쌘��G��(�Y���Y����ޥ���r�WHCy<*��o�|�<a�F��,+�>��~(����[.����N�Dy�Ӵ\ȳ�ۄ޸��`�z`���Y��4���L����93H������&��՚x}P��*�6�}Jz�y���b ��-�c�{)scL��������c!�ɼ��`�@�U?���
��t��O �-�_�I-�"�Б ��;ǹlF;G�