XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170G�jy�,��[��o};�w&���O�e�o�찉��v8Lޏ��X>��z���������r�a��bmL��\��_c������K��q��RP}S؃�S���W	�!�IQ����[Fw �∹4m���u�Q�GW-Jǻ��[�Q�*p��Ǳ�k��$���V�&�Z��-���Sx�s
�vNG���|��!�nR&M/�D�p%<UU ���qP����3]Vǯ���%�c(�"�r�)�*|յ=�r�����rs7�w��g|���Po/���ri��{��r+z4 #��t�k�����OHu�Z�i���C�5��sh�Ͼ�x�$����,#�/�Wi��׽j-"���u���XlxV61EB     400     110�*|�a^���؅a�G&t� (!���#,g��R%Y�>�����^g��|i�a��x���i�C�B�|w���@����� �b���@�,-��
MжW�O�D��{4�VؠDR�d��ܤt�����a�wU:�Cq/�2m��8����D$8�`W��v� G���wOQ#�+D��j��ҿm�
�8��5CV���7@JW!��vFH`�M� "�1�E�&��8`W|�D�#��]��;��i�oF뷞_��)����؆�,�Ǐ�'XlxV61EB     400     120X�i&�;{�F�Y�$���vH c���/h��\eQ�>�_(�^�윢�2�f�d0�A�,����⯔��ni�Z��gHo�E�����F+�]�B������f��qc�飶uO��@�c)�?ĵ^{���!�þ�(���d��n��d��)!E��P�D�(����d0E�ì��r�l����a�)h�z�l_�,�`{��\��=6%�A�-��1�����O�A�XC2!�cj]˽��k�
�	��]�{W��RH�0�& �ƴ��4�XlxV61EB     400     160� .JI �2�Y�6߅3�jU�߂��� �^F"s��v�3P{0�@8�(�DR�04���j؋�&J��G�
�Y��;7��"HW�*���=�	��=2�!J�և~n( /�ɦ�?5$g0!����cq,uE��N�!K�#�F�!T��@Q'6]>�tq5��WfAIYv=$��1+��X��	(��15qq�x<	~�𗤍�w�nUd��]G�4m��>F�����,�b<�]&zV���l��ױ޷�O��+�q����N������9���0N��.���N�k0�Y�`_��5�7�I��e�E�p�x@���g�8ZdGSD�W�����G�]�XlxV61EB     400     180������w��RZ#U2�]`A5�)bPOz='WU&��zE�9CP;7�Y�Ҽ9�+���ܽ���k�W� \�X�b)���Qr���,���N#K���Ƹ�-S@<Ͼ.�6�|�����j��Z�� ,Ͼ��	�>���n��,�Ҿɞk������3��s��er���[J�GqpMb� ^����d�3�8�ⱎ+#t*�zXULMq�����b.�M�ݖ%��{KZ��I�0� �Q\�)���p$�$�U�Jr�Q�%��m�]qv�P_�<)G�>�(�)r��󪀓�n��u9��$�Z@ ��N�'g�q	[��Q�S�\X�"D0��p�L�hb+ ���`�V,�Q{^6�;y\���KB�4?����Y�f��XlxV61EB     400     130Ʀy���؋�aPt�����?��S�3f��bX9V�]�P�١���C�L���JشY澦�'y'N��\:����\���o7�;!�mVA]��ڪ�$=�]����C�QW����Ԣ�K�W��33lF��ݓ�.S�Z�!	v��Ue �C��hO��-���K����R����nN�k�r?����h;�L0�n�k̝Jﱃ�?��Z�r�oyw(��u%q�~	��z����KQ�z-��B���|=�K�.UXH�X��Ywa��6�N�g."1a[�VG9�JK��P��0�*���Z�30XlxV61EB     400     110�K��jւĨ�)�lD,��q�3|��;� e��ŞIT�[pYW�5�#Ұ�j�ݞ��ܳ;S�d6��6V�*X��=��&�Y�	�df�G��Pײ�[��[��f�W�(��ַlh�H*�#������hа���S&���Ny���q�U�H��AS��v�<Ha�P������wE��.��x����<�k<�g�)�y�R�kQYQǥ������DM��{��>�v����jwz����aU,����Ř~ߙ4�?��O��z*XlxV61EB     400      f0�c]������^;T>K�8JP��L�*?s�H�k3ЇF� ��0��������KT� �s��d��6�l�]�.����@~���˲�����چ䟀+ 4�91a�
����$-3�;12�/�ߒ�8�zxS?n�*�R�<���(�d�_Թ
�O����v�#3�����ɍ���c!Dt��̹��<�`ś�dG#�CX͗�:йeM�bk������"W����D�i|��XXlxV61EB     400      c0A�(I�Bi��0\@���^�v�UU�"��r����t������d��ͫIap�؅A�(!�1R	��Y*ϴT��?¡UH�'�^iFv<7�V+����e�_�L���`< ��i�� �GX�׀��%���A�thҪ�y�Ʃ�$"b���mA�?����@b�a<ֵ
8`�K�0��������jރXlxV61EB     400      b0k10ƶ-<q��@���u0(-����+=��J�:��3[%�3Jr����b���i�-,	X��"�4JΤ
]c!���ٮ�	x��C�=���z���κ��{� ��#�����V�5|�yM;�o�$���繄�@xx���b���f��r͖�n�$�@��޾�+Sݓ�M����b+�mXlxV61EB     400     190�轿5��H��btB���8A'��P��q���s޵��5�N�U��
Y/�0����\��n�񧽂��-��(65v����÷5���3Q�ru�P�����=���!��>�-)�w�Ex�u�~W��9V��B�r٤���>r�G	_H;��&�k��t= M�S��=�A�������ҏ����{N��ǃ��⠲Jx������,Thg�Ǟ�n����g�/��9��k��{22�qMP'K���.
��M�U�	U*���o4��G{V��Y��N�P�ӜK���K�W���6!i���!�,� pP�*�s+���}���V�= �ex���9`�dy07_�ў��լ0�'3a�h~A[V��^;�������۴XlxV61EB     400     170�bxذ��w�q��[
�g�Rمq9F�o���	O�V���~�,�� (��X
�q��ʨ�
i�Z@�� +ҕU�U��[©m�)�wh�	��c�A��b\N*,d���ë[#����_��8r6(VoĚ$J����|��Õ��5����
�{��k>N�oLK2Êȏ�Z� ��RS+ػ�[1��i�)�+l#'��$�[��� 		� �;?��y��ǥN��R(�V��a��cOloN��$+�N�*���8
7 26	!l����f��P����e���5�F]����~a�?�u�^;ld)/i��0�v���3��ʘ�S}������η�G���h�I�$ywP_���v��XlxV61EB     400     160��'�Lƕ��zi���Ն>[�UJi���/�v��Χ>�S��=��J��T���ިf��'�pʘ�$�1�c�>��_A����G/��?#�A�C��X�9��q���\���W�����
���	��-���/��<o��i�":�E�(x	3�7�'V5�mf��=�V�5�����uM�b�E���6�i�l/�W�W��Ve�g4��B�k`{��/X��rx�l��L�?� V�'@�cG\)Y"RxVcK���U�kv��5Hh��:�
�W�� =j�ӷȨ>m82s*T�
y�<y�@v���t�a��B=�������úX!Ud�bH��N:�{��o��[�u��XlxV61EB     400     180���@e]�b+n�z�Au���[z��ȩ7N�Q�]`�D_����W`��� ��\�W`Aݜg���y��?�m}aҠ�j�V���3��}G%&2��2j�
��SE��!aC2�ΊZ���H[�bG�"-H�9��,	� ��{�3.o�A���7cZ>-���U�H�G�\�&P�Wz̾!��4���ǔ�_F'Jh�*�RD��H�]@��� Qᴂ(`����1g �s�C܀�Y�ß��C�p-hb�'ȹ/B7q���T�*Cc�+@���g�$W@����E�Y+��2 1�k ^�����pB�;�ws46}�d����Y�검h�!֤��
s5M���i`2�ag��!'�����p��a��STD����&XlxV61EB     400     1a0=�g�|g? 4d!�K���Y�Q�M(�ԃ�5c�H#My���}[_rrg�hM(��)��-(�v�="����x����H&�ծj.���,��6˸#��ф�G��bo�	<�@�cC�:�5������n�}�e�C���-ǲ�P�o�(3���ՍjC��Wd�쾅e4x3`
Ksn�H��2}��Dz�q�s.���+��&�%g���m�������Ǒ��F�	{0�&�J@?�,���n �~�'�f}�4�q�oM��6�U�7�?$?��o�xf�jnH}*$�Ս��������^�e�V$��7��_>��eԲ��e}�[G^��-!�QT�g��Q�p7������q�A�� ��!���;�9E��jy=TWL�p.VTX�`��^�@)o����}�]>XlxV61EB     400      f0�`d!jt=b~DO?��e}�tp�Ao5%	�G 9�F�ӆqzS,�Y�����ܞL��mE	"�T�;�T����K;����٠#j3Xu���� ������U��sP�� ( ����5տt�i��l��N�O���gF]&{����)X�<f�E؎�5���(����,�a�i�q��F���I(�] o^����:�~HTm���^?�h��(�)��u����GTx��;�U[XlxV61EB     400      e0v��J�����@�b���:�Yt�_#E�]��ƕ��2}��^X¤���+la}��]b�F��I�郼��Ӝb�"�� "{ =ՓȈ�p�|��G@��pߡ��{P�5-��th�����
h=����_��y4ժ�Ȑ��"�&�>�`�͸lʢ��(�a�!f��=VX9��5�@�)���)t)i	���oO�v����w2��O��7�~�$���~XlxV61EB     400     100�X�m���5-kR�i�fS�a91u�e�6��Hw��A�� �!�}t�mxL�: ���dڐ�+,_��͙�J>	�Va���@�C�%>}}���Y Tǒ����'M��a�������`�����^�Љ�*P[{\KQ^��;�Ϋ�Q��4\?���zv�X�z�^�j��F�R3��ȿ��YǺ:�M���I�g6�-$xhQ�`l+��C��W�Nn�\��ɂQ13��ՠ��Ѫ��|�M(�fߴ�37s�>XlxV61EB     400     1007Mo��1
�CDS˔�d�*��b�<����*���;�Ɏ���@!a�=aw�����Lu1E��<���ɝK�3��:Eȥy���ܧF���5:n��%�Q���Ը.l�$z�V�[g�6n�ox�Ć����c�#���D4���r��㴫��(ؐn�!�P2�񈢈D��6V���.� ?�,��S>�]ւ׉�Fŧކ�3߾��Y���Ϊe�*?����}��.ka_��Ě0�a^a�V��Z�_-�>`XlxV61EB     400      f0�7��n�>{IMT�s9��i��y�Z�W�p��4<~s��u(ME+���R7���$�Ȳu%9�%��?J�B���?�i�P���kM�Hb.!��l�+�)T���ڳ2�%ꊔg�XM��C<(�q]*��)$=�qJ�E���=��k펠i/Z)H�s����F���?1��s�9<f,o��E�K��2�t>v�I�)����V���ܩJ(�A�y���*�Z�b��8�LCXlxV61EB     400      f07}�F)�w�b����c�05��K�^�`��l"У�4F������!k�%�pvƙ���M��	���[�I[e���|hZ��(�[`y;/�˸���M���R�d��7�`vY*k���&��c�*c�K�ǐ@ؗ�������ױ���/�F�����(S��
zU>�J$����cB��#M�.&�K9!\���y�k*)qC�ǲA��`4���Ϸ���?2ݼ���<;��Q��!XlxV61EB     23e      c0��),��U)/-Gz�����>ј������	5��P��CoE�uo��E(El��7C���j25P��ˉ����d-
$��&5J1�b
Q9錘�#���"�`��]Gkٓ���_^��F�$M�<��n2|@E��vk~��z�(yͦmߥp�T�x�f.�( ��d^�Q6㹜(��㯶�xj�b�