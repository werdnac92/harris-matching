XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     190=9����mf<oi/,|��M���������Խs�BP��H&��q\l	ڇ۬Gt�Ӏna�μ��f[�Gܙ�H(�|�	��E�z��+�����;�*�`~O���ɜ\a�lڏ,t�>��B䒴f�&�]pD)8�����׶�-���gr���^�-��֫�� � ���ҌRg)�q��b�h ��(��Y}�P�/ֹ���X��x���+�dIT f�b����W��u`])����|g����U�۵�0����Q��O^j��<�6J��4T���0{0<�����4#��;Z�Pg��:?(����oX�
�`3r�������E�\�T�����#5KV��.FD>�}Ɣ���B�y����Y����x��ft�e�6";�XlxV61EB     400     140G1^6<��򍃯�jg�=PE�B�|/��%�s0�U~����4H$��5�ǭv�mD -K��ϖ��A��P�����2Zܤ��UR��i0�f ������zŴ0�d���J�"�9?	ćW���Mae�L�����D7<
�?a�cJ���󥂏3o��R����=K��/����M=x+�]�� ��r��y[ܠ���K��2�CdH��~7�v��(��c~t��7�eV�L��*�1�nF0LT�e��x� �|���OR|z� �������X�dU�3�!��#�A@3����4!.�.�W�<�|ĸ��ZY1:j�y�rXlxV61EB     400      e0�W��,�����d����)PR
�8���.�dܟJ`$�%�!��������e � �����C� �:hwF����c�}��0y�a2�#Qn:ʡ&!�8l��+F���x9qe6��أi{���C?�K������eS`y�^��O#jV��KA���Ms'I�'rPj�����Q�lR
v%�6!�O%b���-V���?��A1zw����|V&����o����CDXlxV61EB     400     1b04Q�|_�ζ��^�ԯ*Dj�8Bn�[x�Y�=A�O�,ş0��K���Y�ܟ�
L%l��<��h�Gc���l6Z�n& I��Ӽ���
nc�i�f.�]q�77-@�����ru7ia˙��·�<����bT[���6d�r��o�y����V�2����iTR_<�j��̟%;+�՝��ֿæ���6�]���?gv<O8M�!Qڎ2tN6fS��]�����~ �����`�D���mv�p#����1NnNJ���݈����g�,����^�mS�� ��h����/�eG�B����6Ln��%�E~�R��@���4�/���G�k�uu�"���]�����v�4`�,�]�⪴m&X(���m��o
I۲p��sWy<��n���CO(��?5�ȿ�]� ����!�T�s��]����}XlxV61EB     400     170��p�I[z81ci8�
3��Zc�k�����-o��#��-�t)�L�B�C�#b��B*ū�Np�
�3�)��)xL�SM�J�ei�CW7�5��R������G`���I�.T9s}>��۩6�r��u]+HP�5�G�b(\+�b�zѩ�1#"CJ[�c�����c$u%���j�jsa^kQ*N������fUy-��[������9d߯�)��2؉KH,c�N%���	p0��R�������!۴�FϪ�K�)o�ꛜ՗�j�TM�>7p�X���Ҝ%|�]"n��Z���D8�	�8�J,�~7�]��%JF=�2@���RyRr���2wɢ����)%�;�4=D�����d��6ͧ18��ǧ���XlxV61EB     27c     130�B��t�(�ǕlKA�����"���G]~8��Dcꨱ��[.뱮���8�eC� �a�Slb���>ә��x�+o� ���۲eA�׺���<���7n�p%���]{��/�}́��6A��
߃��NYb�+v%��ι���80���0�*KI$��B�m�}p�����<���VCp�v�|�O�x����1n�:���3�'²�Mt�����x�aT�.1�(%\��]����eRN>B�W�f�[�[�X'a3;�������2���^��\p ,�e�<���_