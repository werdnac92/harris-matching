XlxV61EB     400     140�E�e�?UW�����5�P�x������Z,���[4��$++*�U���"y���A��+�~��N�e�Dt�R��o	C�,��|q�$]�MT�Y��Dͥ�r�N�{ ����x	��-�i;��8tP��P�[2��7b�H9O�V7.�6M�'6�r���w����g���E�D�+�E��h�BYT&�\}�'cgiO(��h�i�,_Zu�n��4�ߖ')��L& I�墰/]݊����,��FR��(�;�R���b�ӎ���s�	���g������g�F�K�W ��֘�6T��WՄ[0�ioK�	;5��Yo`�b^��XlxV61EB     400     170J7Vx1� m�o��������8JA�|�$�m����~�ʬ�{,���-�!���@�{��m�v9U���U��0j��|}��15`N?�_�}&:�@+I�?��CzC�m�Ft\T%nd���?¢� �� ��tXMAc�����U��?�1�j9ruW�q6�y2�����2��ƒUqƦ�P�0K��L��f���5T�{Ϋ>�+^� 4��I�OI�S�8[�u��S���򳃐�j|��b��}�#^����zt(��=�o|2%��6#;�6-�)�/���L�� E:���sj|�\�d}z.����g��;̨pߊy��8�<����ܷ6�4����"���(�����K�3����{|���HsXlxV61EB     400     140A�L��d��2�¿Mj��㧙r�,�)���O�.��/f�/�FFgq,ӭh6�Pd]�P9�����U�K���9�oj��=�=oԖ��CO�
SB���Ȍ`?����z�@kd$��9�eR�)P�~��@�l�z��8&����)�a�m�K��&���h{��15����OW�Q�wtT��U5�R J&�� �)��ñ��Y&ɥ6�с'�T�<b��їZ7�s[���:lߑ�Fp�R��Q�����N��X�ȝ���I���/>�\�" ����-�;t�X�{w૊�~4$3K+��_Er��g�)a�jyXlxV61EB     400     120ן��P�(X��J�i\����]��?�:1\;�%���V�W3MM�c�/��qR��z�c��z"�Ó?���J8�X�m�Jh�,�B:B<#�rgQ;��N��=����K���	�L�@lr�<�Rq��s捔čRK���%�Yx�6�� ���P������B�ܧ1�:ًa�D;@�UlC��"g��}u�Z=ق!�<�V��]_~�����躝!І(!w!P�~E���c��V��� 2����N��gY��B�pf���0�J>k�b�UG�	��g�@�XlxV61EB     400     100�sG&�?�$�p�	7�.AZ)�n���������z�#�~3��yŖ�UA�M ��dʬv9ɹ]!��ڟ'�S۹�(���>�����4_&�.��h*�?�3�/er�!7&�E�/���bL;�Jcܾ�x�?��X��/D	Z��qDVU����
�� ԣq�a�	�~�&��خ����8ߘ�m%�3S]xp\��.���w����X-���9E��6_�V�pP����T��˷^w�ud��U�XlxV61EB     123      c0J��#sQ��A#��:x�Q���~2�DI�Z�2<�"4�甦�*4l�����v8%����i;!��
��h�C�0�,�Ź��!�W���>!����5��D��s�h9�.� cW>�ZB�1_SĊהhJB�� �Xk2�k�~���q��[���ݪ����C�h:�B�Y4�nx���[��j���B|_