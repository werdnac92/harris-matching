XlxV61EB     400     130{�0� �gA�b�DA��vB�~���	)����@� �˷;i��U�\���c�O���F�:�)^���Ү6:�L;��k�J�r+��ff���v	�BI*&T�Qx�b��pL��7xg�cQ[p��[zj� }ɶ�ඝ����G(�q6�{3|�:�W�jۙ^c�ְ�Z`wٟ�i�R
/����)�pXç���ſ���X��-I�}�!it�V����?�����Ҙ�6��(#bl���"0?G����_�g[�
�m�C<&3�7�.:卥��G/eNF��&�XlxV61EB     400     170���H��S@ڐ��|��49ڏ��6�+y�X������3'4Bj���o%�EjKd�tB1��)$�b���5Ϳ	#�l�6�����i�$��ɒ���2
��P�2��h.�sR�e�j��tl~՟�Eyo�9j@�ː2��V��|�"�\���\��|��	M�~���)�J�9�o5[�FY���=��#N��Kue>>�Ht��q��0�C�skl�Z�$i�J0��3a�3Q����S}��".m��՞��d�м�qb'���s����y��O3S��O�U�:���|LMW���a+C!�P��_�l�{��݀�m�� X�!Q2N���5�r�����q��G��CC�\��f��1�K9�܇������XlxV61EB     400     1c0�Ho=*A����K�^���;r��P"�T z�#��P�Yw�3��i��i�k�-��HMW�W×��3�[ٳ��V��OPz�^G�\'���qk��ދO�V8�H\ifhK�z����g0CQ�`��������tlх9j�����@/�����!���H+,��(!J�TJ����~̯p`3�H?��5�Ve9�Bw��.�����v�V�v�2�@�m��,(Caw�*@>��ɇ�`�_^ñ���6��|${ �\� ��,ȲY��,����Hu����$�� �d	��A�E���Ět���Ras~��o�Xva2�[��[��݅+��B<�J򲯜�6���w�a�&ݍ��(q����G��@��me����0��W#��j�A����P Y�ө �o��4-��_��պ�dPO5Я���N���:��5_XlxV61EB     400     160�|�9p
��2�	k���?��{YQL�e�y�ş�R_�V6�b�ɀ��nqؒG���#X٧&��е-�����	�c-��4�Gd�q�80����P^�o2����՜`ݯ���r�(e�=��,V����jV��4.co٭�����fʐUڍ�������Vt9-*;p�����8�+gŴ���sJ'}��i��e I�(�9��������?���B�M{��B�)8Ì����%E԰X��@ò����<�'����.���ܬ3������c���h�:���������<�D��kU�jr^�,��1$�\����<#�u�{�~�Xo`��nɒ�7�j/��u�Ԝ��XlxV61EB     121      a0o�?/"��P|��n���x�O$s���9��|�&+���AH&U.[.��r����ڔ�I��6X����T�+�7_F��~�W��D&��Ig��@K�ӆ�)\�BZ����>c��R񲀁m,�i�	�e��gg����nR��`�.&uCgg%��